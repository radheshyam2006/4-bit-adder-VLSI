.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u

vdd vdd gnd DC 1.8

.subckt nmos d g s b W='N'
.param width_N={W}
M1 d g s b CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends nmos

.subckt pmos d g s b W='P'
.param width_P={W}
M1 d g s b CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends pmos

.subckt inv out in vdd gnd N='a'
.param width_N={N}
.param width_P={2*width_N}
M1      out       in      gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      out       in      vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

.subckt xor out a b clk vdd gnd
Xabar abar a vdd gnd inv N='10*LAMBDA'
Xbbar bbar b vdd gnd inv N='10*LAMBDA'

X1 n12 abar vdd vdd pmos W='20*LAMBDA'
X2 n23 bbar n12 n12 pmos W='20*LAMBDA'
X3 n67 a vdd vdd pmos W='20*LAMBDA'
X4 n23 b n67 n67 pmos W='20*LAMBDA'
X5 n34 clk n23 n23 pmos W='20*LAMBDA'
X6 n34 abar n45 n45 nmos W='10*LAMBDA'
X7 n45 b gnd gnd nmos W='10*LAMBDA'
X8 n34 a n89 n89 nmos W='10*LAMBDA'
X9 n89 bbar gnd gnd nmos W='10*LAMBDA'

X10 m67 n34 vdd vdd pmos W='20*LAMBDA'
X11 m78 clk m67 m67 pmos W='20*LAMBDA'
X12 m78 n34 gnd gnd nmos W='10*LAMBDA'

X13 m910 m78 vdd vdd pmos W='20*LAMBDA'
X14 m910 clk m1011 m1011 nmos W='10*LAMBDA'
X15 m1011 m78 gnd gnd nmos W='10*LAMBDA'

X16 out m910 vdd vdd pmos W='20*LAMBDA'
X17 out clk m1314 m1314 nmos W='10*LAMBDA'
X18 m1314 m910 gnd gnd nmos W='10*LAMBDA'
.ends xor

V1 clk gnd pulse(0 1.8 80n 0 0 40n 80n)
V2 a gnd pulse(0 1.8 10n 0 0 160n 320n)
V3 b gnd pulse(0 1.8 15n 0 0 320n 640n)

Xxor out a b clk vdd gnd xor

.tran 0.1n 640ns
.control
run
set hcopypscolor = 1
set color0 = white
set color1 = blue
plot v(clk) v(a)+6 v(b)+4 v(out)+2
.endc
