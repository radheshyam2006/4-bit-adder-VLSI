magic
tech scmos
timestamp 1732004181
<< nwell >>
rect -729 969 -696 1016
rect -665 973 -633 1011
rect -249 872 -221 906
rect -552 775 -519 822
rect -500 781 -434 823
rect -219 782 -191 836
rect -723 685 -690 732
rect -659 689 -627 727
rect -235 723 -207 757
rect -182 754 -154 778
rect -253 634 -225 668
rect -548 533 -515 580
rect -496 539 -430 581
rect -223 544 -195 598
rect -28 541 5 588
rect 24 547 90 589
rect -239 485 -211 519
rect -186 516 -158 540
rect -711 429 -678 476
rect -647 433 -615 471
rect -248 407 -220 441
rect -536 299 -503 346
rect -484 305 -418 347
rect -218 317 -190 371
rect -24 319 9 366
rect 28 325 94 367
rect -234 258 -206 292
rect -181 289 -153 313
rect -246 184 -218 218
rect -688 54 -655 101
rect -624 58 -592 96
rect -529 83 -496 130
rect -477 89 -411 131
rect -216 94 -188 148
rect -17 106 16 153
rect 35 112 101 154
rect -232 35 -204 69
rect -179 66 -151 90
rect -8 -67 25 -20
rect 44 -61 110 -19
<< ntransistor >>
rect -713 951 -711 961
rect -651 942 -649 952
rect -660 890 -658 900
rect -237 852 -235 862
rect -536 757 -534 767
rect -328 782 -326 823
rect -321 782 -319 823
rect -295 783 -293 823
rect -268 783 -266 823
rect -245 783 -243 823
rect -487 754 -485 764
rect -453 754 -451 764
rect -342 705 -340 745
rect -318 705 -316 745
rect -297 705 -295 745
rect -280 705 -278 745
rect -262 706 -260 746
rect -223 703 -221 713
rect -707 667 -705 677
rect -645 658 -643 668
rect -654 606 -652 616
rect -241 614 -239 624
rect -532 515 -530 525
rect -315 544 -313 585
rect -308 544 -306 585
rect -282 545 -280 585
rect -255 545 -253 585
rect -483 512 -481 522
rect -449 512 -447 522
rect -329 467 -327 507
rect -305 467 -303 507
rect -284 467 -282 507
rect -267 467 -265 507
rect -12 523 -10 533
rect 37 520 39 530
rect 71 520 73 530
rect -227 465 -225 475
rect -695 411 -693 421
rect -633 402 -631 412
rect -236 387 -234 397
rect -642 350 -640 360
rect -520 281 -518 291
rect -283 317 -281 358
rect -276 317 -274 358
rect -250 318 -248 358
rect -8 301 -6 311
rect 41 298 43 308
rect 75 298 77 308
rect -471 278 -469 288
rect -437 278 -435 288
rect -297 240 -295 280
rect -273 240 -271 280
rect -252 240 -250 280
rect -222 238 -220 248
rect -234 164 -232 174
rect -513 65 -511 75
rect -262 94 -260 135
rect -255 94 -253 135
rect -1 88 1 98
rect 48 85 50 95
rect 82 85 84 95
rect -464 62 -462 72
rect -430 62 -428 72
rect -672 36 -670 46
rect -610 27 -608 37
rect -276 17 -274 57
rect -252 17 -250 57
rect -220 15 -218 25
rect -619 -25 -617 -15
rect 8 -85 10 -75
rect 57 -88 59 -78
rect 91 -88 93 -78
<< ptransistor >>
rect -713 981 -711 1001
rect -651 984 -649 1004
rect -237 880 -235 900
rect -536 787 -534 807
rect -487 795 -485 815
rect -453 795 -451 815
rect -207 790 -205 830
rect -170 762 -168 772
rect -707 697 -705 717
rect -645 700 -643 720
rect -223 731 -221 751
rect -241 642 -239 662
rect -532 545 -530 565
rect -483 553 -481 573
rect -449 553 -447 573
rect -211 552 -209 592
rect -12 553 -10 573
rect 37 561 39 581
rect 71 561 73 581
rect -174 524 -172 534
rect -227 493 -225 513
rect -695 441 -693 461
rect -633 444 -631 464
rect -236 415 -234 435
rect -520 311 -518 331
rect -471 319 -469 339
rect -437 319 -435 339
rect -206 325 -204 365
rect -8 331 -6 351
rect 41 339 43 359
rect 75 339 77 359
rect -169 297 -167 307
rect -222 266 -220 286
rect -234 192 -232 212
rect -513 95 -511 115
rect -464 103 -462 123
rect -430 103 -428 123
rect -672 66 -670 86
rect -610 69 -608 89
rect -204 102 -202 142
rect -1 118 1 138
rect 48 126 50 146
rect 82 126 84 146
rect -167 74 -165 84
rect -220 43 -218 63
rect 8 -55 10 -35
rect 57 -47 59 -27
rect 91 -47 93 -27
<< ndiffusion >>
rect -714 951 -713 961
rect -711 951 -710 961
rect -652 942 -651 952
rect -649 942 -648 952
rect -661 890 -660 900
rect -658 890 -657 900
rect -238 852 -237 862
rect -235 852 -234 862
rect -537 757 -536 767
rect -534 757 -533 767
rect -329 782 -328 823
rect -326 782 -321 823
rect -319 782 -318 823
rect -296 783 -295 823
rect -293 783 -292 823
rect -269 783 -268 823
rect -266 783 -265 823
rect -246 783 -245 823
rect -243 783 -242 823
rect -488 754 -487 764
rect -485 754 -484 764
rect -454 754 -453 764
rect -451 754 -450 764
rect -343 705 -342 745
rect -340 705 -339 745
rect -319 705 -318 745
rect -316 705 -315 745
rect -298 705 -297 745
rect -295 705 -294 745
rect -281 705 -280 745
rect -278 705 -277 745
rect -263 706 -262 746
rect -260 706 -259 746
rect -224 703 -223 713
rect -221 703 -220 713
rect -708 667 -707 677
rect -705 667 -704 677
rect -646 658 -645 668
rect -643 658 -642 668
rect -655 606 -654 616
rect -652 606 -651 616
rect -242 614 -241 624
rect -239 614 -238 624
rect -533 515 -532 525
rect -530 515 -529 525
rect -316 544 -315 585
rect -313 544 -308 585
rect -306 544 -305 585
rect -283 545 -282 585
rect -280 545 -279 585
rect -256 545 -255 585
rect -253 545 -252 585
rect -484 512 -483 522
rect -481 512 -480 522
rect -450 512 -449 522
rect -447 512 -446 522
rect -330 467 -329 507
rect -327 467 -326 507
rect -306 467 -305 507
rect -303 467 -302 507
rect -285 467 -284 507
rect -282 467 -281 507
rect -268 467 -267 507
rect -265 467 -264 507
rect -13 523 -12 533
rect -10 523 -9 533
rect 36 520 37 530
rect 39 520 40 530
rect 70 520 71 530
rect 73 520 74 530
rect -228 465 -227 475
rect -225 465 -224 475
rect -696 411 -695 421
rect -693 411 -692 421
rect -634 402 -633 412
rect -631 402 -630 412
rect -237 387 -236 397
rect -234 387 -233 397
rect -643 350 -642 360
rect -640 350 -639 360
rect -521 281 -520 291
rect -518 281 -517 291
rect -284 317 -283 358
rect -281 317 -276 358
rect -274 317 -273 358
rect -251 318 -250 358
rect -248 318 -247 358
rect -9 301 -8 311
rect -6 301 -5 311
rect 40 298 41 308
rect 43 298 44 308
rect 74 298 75 308
rect 77 298 78 308
rect -472 278 -471 288
rect -469 278 -468 288
rect -438 278 -437 288
rect -435 278 -434 288
rect -298 240 -297 280
rect -295 240 -294 280
rect -274 240 -273 280
rect -271 240 -270 280
rect -253 240 -252 280
rect -250 240 -249 280
rect -223 238 -222 248
rect -220 238 -219 248
rect -235 164 -234 174
rect -232 164 -231 174
rect -514 65 -513 75
rect -511 65 -510 75
rect -263 94 -262 135
rect -260 94 -255 135
rect -253 94 -252 135
rect -2 88 -1 98
rect 1 88 2 98
rect 47 85 48 95
rect 50 85 51 95
rect 81 85 82 95
rect 84 85 85 95
rect -465 62 -464 72
rect -462 62 -461 72
rect -431 62 -430 72
rect -428 62 -427 72
rect -673 36 -672 46
rect -670 36 -669 46
rect -611 27 -610 37
rect -608 27 -607 37
rect -277 17 -276 57
rect -274 17 -273 57
rect -253 17 -252 57
rect -250 17 -249 57
rect -221 15 -220 25
rect -218 15 -217 25
rect -620 -25 -619 -15
rect -617 -25 -616 -15
rect 7 -85 8 -75
rect 10 -85 11 -75
rect 56 -88 57 -78
rect 59 -88 60 -78
rect 90 -88 91 -78
rect 93 -88 94 -78
<< pdiffusion >>
rect -714 981 -713 1001
rect -711 981 -710 1001
rect -652 984 -651 1004
rect -649 984 -648 1004
rect -238 880 -237 900
rect -235 880 -234 900
rect -537 787 -536 807
rect -534 787 -533 807
rect -488 795 -487 815
rect -485 795 -484 815
rect -454 795 -453 815
rect -451 795 -450 815
rect -208 790 -207 830
rect -205 790 -204 830
rect -171 762 -170 772
rect -168 762 -167 772
rect -708 697 -707 717
rect -705 697 -704 717
rect -646 700 -645 720
rect -643 700 -642 720
rect -224 731 -223 751
rect -221 731 -220 751
rect -242 642 -241 662
rect -239 642 -238 662
rect -533 545 -532 565
rect -530 545 -529 565
rect -484 553 -483 573
rect -481 553 -480 573
rect -450 553 -449 573
rect -447 553 -446 573
rect -212 552 -211 592
rect -209 552 -208 592
rect -13 553 -12 573
rect -10 553 -9 573
rect 36 561 37 581
rect 39 561 40 581
rect 70 561 71 581
rect 73 561 74 581
rect -175 524 -174 534
rect -172 524 -171 534
rect -228 493 -227 513
rect -225 493 -224 513
rect -696 441 -695 461
rect -693 441 -692 461
rect -634 444 -633 464
rect -631 444 -630 464
rect -237 415 -236 435
rect -234 415 -233 435
rect -521 311 -520 331
rect -518 311 -517 331
rect -472 319 -471 339
rect -469 319 -468 339
rect -438 319 -437 339
rect -435 319 -434 339
rect -207 325 -206 365
rect -204 325 -203 365
rect -9 331 -8 351
rect -6 331 -5 351
rect 40 339 41 359
rect 43 339 44 359
rect 74 339 75 359
rect 77 339 78 359
rect -170 297 -169 307
rect -167 297 -166 307
rect -223 266 -222 286
rect -220 266 -219 286
rect -235 192 -234 212
rect -232 192 -231 212
rect -514 95 -513 115
rect -511 95 -510 115
rect -465 103 -464 123
rect -462 103 -461 123
rect -431 103 -430 123
rect -428 103 -427 123
rect -673 66 -672 86
rect -670 66 -669 86
rect -611 69 -610 89
rect -608 69 -607 89
rect -205 102 -204 142
rect -202 102 -201 142
rect -2 118 -1 138
rect 1 118 2 138
rect 47 126 48 146
rect 50 126 51 146
rect 81 126 82 146
rect 84 126 85 146
rect -168 74 -167 84
rect -165 74 -164 84
rect -221 43 -220 63
rect -218 43 -217 63
rect 7 -55 8 -35
rect 10 -55 11 -35
rect 56 -47 57 -27
rect 59 -47 60 -27
rect 90 -47 91 -27
rect 93 -47 94 -27
<< ndcontact >>
rect -718 951 -714 961
rect -710 951 -706 961
rect -656 942 -652 952
rect -648 942 -644 952
rect -665 890 -661 900
rect -657 890 -653 900
rect -242 852 -238 862
rect -234 852 -230 862
rect -541 757 -537 767
rect -533 757 -529 767
rect -333 782 -329 823
rect -318 782 -313 823
rect -300 783 -296 823
rect -292 783 -288 823
rect -273 783 -269 823
rect -265 783 -261 823
rect -250 783 -246 823
rect -242 783 -238 823
rect -492 754 -488 764
rect -484 754 -480 764
rect -458 754 -454 764
rect -450 754 -446 764
rect -347 705 -343 745
rect -339 705 -335 745
rect -323 705 -319 745
rect -315 705 -311 745
rect -302 705 -298 745
rect -294 705 -290 745
rect -285 705 -281 745
rect -277 705 -273 745
rect -267 706 -263 746
rect -259 706 -255 746
rect -228 703 -224 713
rect -220 703 -216 713
rect -712 667 -708 677
rect -704 667 -700 677
rect -650 658 -646 668
rect -642 658 -638 668
rect -659 606 -655 616
rect -651 606 -647 616
rect -246 614 -242 624
rect -238 614 -234 624
rect -537 515 -533 525
rect -529 515 -525 525
rect -320 544 -316 585
rect -305 544 -300 585
rect -287 545 -283 585
rect -279 545 -275 585
rect -260 545 -256 585
rect -252 545 -248 585
rect -488 512 -484 522
rect -480 512 -476 522
rect -454 512 -450 522
rect -446 512 -442 522
rect -334 467 -330 507
rect -326 467 -322 507
rect -310 467 -306 507
rect -302 467 -298 507
rect -289 467 -285 507
rect -281 467 -277 507
rect -272 467 -268 507
rect -264 467 -260 507
rect -17 523 -13 533
rect -9 523 -5 533
rect 32 520 36 530
rect 40 520 44 530
rect 66 520 70 530
rect 74 520 78 530
rect -232 465 -228 475
rect -224 465 -220 475
rect -700 411 -696 421
rect -692 411 -688 421
rect -638 402 -634 412
rect -630 402 -626 412
rect -241 387 -237 397
rect -233 387 -229 397
rect -647 350 -643 360
rect -639 350 -635 360
rect -525 281 -521 291
rect -517 281 -513 291
rect -288 317 -284 358
rect -273 317 -268 358
rect -255 318 -251 358
rect -247 318 -243 358
rect -13 301 -9 311
rect -5 301 -1 311
rect 36 298 40 308
rect 44 298 48 308
rect 70 298 74 308
rect 78 298 82 308
rect -476 278 -472 288
rect -468 278 -464 288
rect -442 278 -438 288
rect -434 278 -430 288
rect -302 240 -298 280
rect -294 240 -290 280
rect -278 240 -274 280
rect -270 240 -266 280
rect -257 240 -253 280
rect -249 240 -245 280
rect -227 238 -223 248
rect -219 238 -215 248
rect -239 164 -235 174
rect -231 164 -227 174
rect -518 65 -514 75
rect -510 65 -506 75
rect -267 94 -263 135
rect -252 94 -247 135
rect -6 88 -2 98
rect 2 88 6 98
rect 43 85 47 95
rect 51 85 55 95
rect 77 85 81 95
rect 85 85 89 95
rect -469 62 -465 72
rect -461 62 -457 72
rect -435 62 -431 72
rect -427 62 -423 72
rect -677 36 -673 46
rect -669 36 -665 46
rect -615 27 -611 37
rect -607 27 -603 37
rect -281 17 -277 57
rect -273 17 -269 57
rect -257 17 -253 57
rect -249 17 -245 57
rect -225 15 -221 25
rect -217 15 -213 25
rect -624 -25 -620 -15
rect -616 -25 -612 -15
rect 3 -85 7 -75
rect 11 -85 15 -75
rect 52 -88 56 -78
rect 60 -88 64 -78
rect 86 -88 90 -78
rect 94 -88 98 -78
<< pdcontact >>
rect -718 981 -714 1001
rect -710 981 -706 1001
rect -656 984 -652 1004
rect -648 984 -644 1004
rect -242 880 -238 900
rect -234 880 -230 900
rect -541 787 -537 807
rect -533 787 -529 807
rect -492 795 -488 815
rect -484 795 -480 815
rect -458 795 -454 815
rect -450 795 -446 815
rect -212 790 -208 830
rect -204 790 -200 830
rect -175 762 -171 772
rect -167 762 -163 772
rect -712 697 -708 717
rect -704 697 -700 717
rect -650 700 -646 720
rect -642 700 -638 720
rect -228 731 -224 751
rect -220 731 -216 751
rect -246 642 -242 662
rect -238 642 -234 662
rect -537 545 -533 565
rect -529 545 -525 565
rect -488 553 -484 573
rect -480 553 -476 573
rect -454 553 -450 573
rect -446 553 -442 573
rect -216 552 -212 592
rect -208 552 -204 592
rect -17 553 -13 573
rect -9 553 -5 573
rect 32 561 36 581
rect 40 561 44 581
rect 66 561 70 581
rect 74 561 78 581
rect -179 524 -175 534
rect -171 524 -167 534
rect -232 493 -228 513
rect -224 493 -220 513
rect -700 441 -696 461
rect -692 441 -688 461
rect -638 444 -634 464
rect -630 444 -626 464
rect -241 415 -237 435
rect -233 415 -229 435
rect -525 311 -521 331
rect -517 311 -513 331
rect -476 319 -472 339
rect -468 319 -464 339
rect -442 319 -438 339
rect -434 319 -430 339
rect -211 325 -207 365
rect -203 325 -199 365
rect -13 331 -9 351
rect -5 331 -1 351
rect 36 339 40 359
rect 44 339 48 359
rect 70 339 74 359
rect 78 339 82 359
rect -174 297 -170 307
rect -166 297 -162 307
rect -227 266 -223 286
rect -219 266 -215 286
rect -239 192 -235 212
rect -231 192 -227 212
rect -518 95 -514 115
rect -510 95 -506 115
rect -469 103 -465 123
rect -461 103 -457 123
rect -435 103 -431 123
rect -427 103 -423 123
rect -677 66 -673 86
rect -669 66 -665 86
rect -615 69 -611 89
rect -607 69 -603 89
rect -209 102 -205 142
rect -201 102 -197 142
rect -6 118 -2 138
rect 2 118 6 138
rect 43 126 47 146
rect 51 126 55 146
rect 77 126 81 146
rect 85 126 89 146
rect -172 74 -168 84
rect -164 74 -160 84
rect -225 43 -221 63
rect -217 43 -213 63
rect 3 -55 7 -35
rect 11 -55 15 -35
rect 52 -47 56 -27
rect 60 -47 64 -27
rect 86 -47 90 -27
rect 94 -47 98 -27
<< polysilicon >>
rect -713 1001 -711 1010
rect -651 1004 -649 1014
rect -713 961 -711 981
rect -651 969 -649 984
rect -651 952 -649 957
rect -713 948 -711 951
rect -651 937 -649 942
rect -660 900 -658 921
rect -237 900 -235 903
rect -660 883 -658 890
rect -237 862 -235 880
rect -237 849 -235 852
rect -207 830 -205 833
rect -328 823 -326 830
rect -321 823 -319 830
rect -295 823 -293 830
rect -268 823 -266 830
rect -245 823 -243 830
rect -536 807 -534 816
rect -487 815 -485 822
rect -453 815 -451 819
rect -536 767 -534 787
rect -487 780 -485 795
rect -487 764 -485 767
rect -453 764 -451 795
rect -328 779 -326 782
rect -321 779 -319 782
rect -295 779 -293 783
rect -268 779 -266 783
rect -245 779 -243 783
rect -207 775 -205 790
rect -170 772 -168 775
rect -536 754 -534 757
rect -487 735 -485 754
rect -453 751 -451 754
rect -342 745 -340 752
rect -318 745 -316 752
rect -297 745 -295 752
rect -280 745 -278 752
rect -262 746 -260 753
rect -223 751 -221 754
rect -707 717 -705 726
rect -645 720 -643 730
rect -170 747 -168 762
rect -223 713 -221 731
rect -342 701 -340 705
rect -318 701 -316 705
rect -297 701 -295 705
rect -280 701 -278 705
rect -262 702 -260 706
rect -223 700 -221 703
rect -707 677 -705 697
rect -645 685 -643 700
rect -645 668 -643 673
rect -707 664 -705 667
rect -241 662 -239 665
rect -645 653 -643 658
rect -654 616 -652 637
rect -241 624 -239 642
rect -241 611 -239 614
rect -654 599 -652 606
rect -211 592 -209 595
rect -315 585 -313 592
rect -308 585 -306 592
rect -282 585 -280 592
rect -255 585 -253 592
rect -532 565 -530 574
rect -483 573 -481 580
rect -449 573 -447 577
rect -532 525 -530 545
rect -483 538 -481 553
rect -483 522 -481 525
rect -449 522 -447 553
rect -12 573 -10 582
rect 37 581 39 588
rect 71 581 73 585
rect -315 541 -313 544
rect -308 541 -306 544
rect -282 541 -280 545
rect -255 541 -253 545
rect -211 537 -209 552
rect -174 534 -172 537
rect -12 533 -10 553
rect 37 546 39 561
rect -532 512 -530 515
rect -483 493 -481 512
rect -449 509 -447 512
rect -329 507 -327 514
rect -305 507 -303 514
rect -284 507 -282 514
rect -267 507 -265 514
rect -227 513 -225 516
rect -695 461 -693 470
rect -633 464 -631 474
rect -174 509 -172 524
rect 37 530 39 533
rect 71 530 73 561
rect -12 520 -10 523
rect 37 501 39 520
rect 71 517 73 520
rect -227 475 -225 493
rect -329 463 -327 467
rect -305 463 -303 467
rect -284 463 -282 467
rect -267 463 -265 467
rect -227 462 -225 465
rect -695 421 -693 441
rect -633 429 -631 444
rect -236 435 -234 438
rect -633 412 -631 417
rect -695 408 -693 411
rect -633 397 -631 402
rect -236 397 -234 415
rect -236 384 -234 387
rect -642 360 -640 381
rect -206 365 -204 368
rect -283 358 -281 365
rect -276 358 -274 365
rect -250 358 -248 365
rect -642 343 -640 350
rect -520 331 -518 340
rect -471 339 -469 346
rect -437 339 -435 343
rect -520 291 -518 311
rect -471 304 -469 319
rect -471 288 -469 291
rect -437 288 -435 319
rect -8 351 -6 360
rect 41 359 43 366
rect 75 359 77 363
rect -283 314 -281 317
rect -276 314 -274 317
rect -250 314 -248 318
rect -206 310 -204 325
rect -8 311 -6 331
rect 41 324 43 339
rect -169 307 -167 310
rect 41 308 43 311
rect 75 308 77 339
rect -8 298 -6 301
rect -520 278 -518 281
rect -297 280 -295 287
rect -273 280 -271 287
rect -252 280 -250 287
rect -222 286 -220 289
rect -471 259 -469 278
rect -437 275 -435 278
rect -169 282 -167 297
rect 41 279 43 298
rect 75 295 77 298
rect -222 248 -220 266
rect -297 236 -295 240
rect -273 236 -271 240
rect -252 236 -250 240
rect -222 235 -220 238
rect -234 212 -232 215
rect -234 174 -232 192
rect -234 161 -232 164
rect -204 142 -202 145
rect -262 135 -260 142
rect -255 135 -253 142
rect -513 115 -511 124
rect -464 123 -462 130
rect -430 123 -428 127
rect -672 86 -670 95
rect -610 89 -608 99
rect -513 75 -511 95
rect -464 88 -462 103
rect -672 46 -670 66
rect -610 54 -608 69
rect -464 72 -462 75
rect -430 72 -428 103
rect -1 138 1 147
rect 48 146 50 153
rect 82 146 84 150
rect -262 91 -260 94
rect -255 91 -253 94
rect -204 87 -202 102
rect -1 98 1 118
rect 48 111 50 126
rect 48 95 50 98
rect 82 95 84 126
rect -167 84 -165 87
rect -1 85 1 88
rect -513 62 -511 65
rect -464 43 -462 62
rect -430 59 -428 62
rect -276 57 -274 64
rect -252 57 -250 64
rect -220 63 -218 66
rect -610 37 -608 42
rect -672 33 -670 36
rect -610 22 -608 27
rect -167 59 -165 74
rect 48 66 50 85
rect 82 82 84 85
rect -220 25 -218 43
rect -276 13 -274 17
rect -252 13 -250 17
rect -220 12 -218 15
rect -619 -15 -617 6
rect -619 -32 -617 -25
rect 8 -35 10 -26
rect 57 -27 59 -20
rect 91 -27 93 -23
rect 8 -75 10 -55
rect 57 -62 59 -47
rect 57 -78 59 -75
rect 91 -78 93 -47
rect 8 -88 10 -85
rect 57 -107 59 -88
rect 91 -91 93 -88
<< polycontact >>
rect -655 1014 -649 1021
rect -717 964 -713 968
rect -655 930 -649 937
rect -662 921 -658 925
rect -241 866 -237 870
rect -332 826 -328 830
rect -319 826 -315 830
rect -299 826 -295 830
rect -272 826 -268 830
rect -249 826 -245 830
rect -485 818 -481 822
rect -540 770 -536 774
rect -457 771 -453 775
rect -211 775 -207 779
rect -649 730 -643 737
rect -346 748 -342 752
rect -322 748 -318 752
rect -301 748 -297 752
rect -284 748 -280 752
rect -266 749 -262 753
rect -485 735 -480 740
rect -174 747 -170 751
rect -227 717 -223 721
rect -711 680 -707 684
rect -649 646 -643 653
rect -656 637 -652 641
rect -245 628 -241 632
rect -319 588 -315 592
rect -306 588 -302 592
rect -286 588 -282 592
rect -259 588 -255 592
rect -481 576 -477 580
rect -536 528 -532 532
rect -453 529 -449 533
rect 39 584 43 588
rect -215 537 -211 541
rect -16 536 -12 540
rect 67 537 71 541
rect -333 510 -329 514
rect -309 510 -305 514
rect -288 510 -284 514
rect -271 510 -267 514
rect -481 493 -476 498
rect -637 474 -631 481
rect -178 509 -174 513
rect 39 501 44 506
rect -231 479 -227 483
rect -699 424 -695 428
rect -240 401 -236 405
rect -637 390 -631 397
rect -644 381 -640 385
rect -287 361 -283 365
rect -274 361 -270 365
rect -254 361 -250 365
rect -469 342 -465 346
rect -524 294 -520 298
rect -441 295 -437 299
rect 43 362 47 366
rect -210 310 -206 314
rect -12 314 -8 318
rect 71 315 75 319
rect -301 283 -297 287
rect -277 283 -273 287
rect -256 283 -252 287
rect -469 259 -464 264
rect -173 282 -169 286
rect 43 279 48 284
rect -226 252 -222 256
rect -238 178 -234 182
rect -266 138 -262 142
rect -253 138 -249 142
rect -462 126 -458 130
rect -614 99 -608 106
rect -517 78 -513 82
rect -434 79 -430 83
rect -676 49 -672 53
rect 50 149 54 153
rect -208 87 -204 91
rect -5 101 -1 105
rect 78 102 82 106
rect -280 60 -276 64
rect -256 60 -252 64
rect -462 43 -457 48
rect -614 15 -608 22
rect -171 59 -167 63
rect 50 66 55 71
rect -224 29 -220 33
rect -621 6 -617 10
rect 59 -24 63 -20
rect 4 -72 8 -68
rect 87 -71 91 -67
rect 59 -107 64 -102
<< metal1 >>
rect -754 1026 -680 1031
rect -754 899 -748 1026
rect -729 1016 -696 1023
rect -684 1021 -680 1026
rect -718 1001 -714 1016
rect -684 1014 -655 1021
rect -742 968 -737 971
rect -742 964 -717 968
rect -710 967 -706 981
rect -684 971 -677 1014
rect -687 967 -677 971
rect -742 963 -734 964
rect -710 963 -683 967
rect -656 965 -652 984
rect -742 917 -737 963
rect -710 961 -706 963
rect -673 959 -652 965
rect -656 952 -652 959
rect -718 946 -714 951
rect -729 939 -693 946
rect -648 966 -644 984
rect -648 960 -613 966
rect -648 952 -644 960
rect -681 930 -655 937
rect -681 917 -674 930
rect -742 911 -674 917
rect -670 921 -662 925
rect -670 907 -667 921
rect -619 917 -613 960
rect -673 903 -667 907
rect -657 911 -613 917
rect -673 899 -670 903
rect -657 900 -653 911
rect -249 906 -221 909
rect -754 895 -670 899
rect -242 900 -239 906
rect -665 877 -661 890
rect -677 872 -641 877
rect -233 870 -230 880
rect -249 866 -241 870
rect -233 867 -221 870
rect -233 862 -230 867
rect -509 845 -502 854
rect -475 836 -468 852
rect -242 844 -239 852
rect -249 841 -239 844
rect -227 838 -224 840
rect -567 832 -468 836
rect -567 774 -558 832
rect -552 822 -509 829
rect -475 822 -468 832
rect -335 826 -332 830
rect -315 826 -309 830
rect -302 826 -299 830
rect -275 826 -272 830
rect -252 826 -249 830
rect -242 829 -238 830
rect -242 825 -231 829
rect -242 823 -238 825
rect -541 807 -537 822
rect -481 818 -454 822
rect -458 815 -454 818
rect -567 770 -540 774
rect -533 773 -529 787
rect -492 776 -488 795
rect -533 769 -506 773
rect -533 767 -529 769
rect -541 752 -537 757
rect -748 742 -674 747
rect -552 745 -516 752
rect -748 615 -742 742
rect -723 732 -690 739
rect -678 737 -674 742
rect -712 717 -708 732
rect -678 730 -649 737
rect -511 731 -506 769
rect -492 764 -488 770
rect -492 748 -488 754
rect -484 764 -480 795
rect -450 776 -446 795
rect -464 771 -457 775
rect -450 770 -427 776
rect -333 773 -329 782
rect -318 781 -313 782
rect -300 781 -296 783
rect -318 776 -296 781
rect -292 781 -288 783
rect -273 781 -269 783
rect -292 776 -269 781
rect -265 781 -261 783
rect -250 781 -246 783
rect -265 776 -246 781
rect -450 764 -446 770
rect -338 769 -320 773
rect -463 758 -458 764
rect -484 747 -480 754
rect -450 747 -446 754
rect -349 748 -346 752
rect -484 743 -446 747
rect -339 745 -335 754
rect -480 735 -476 740
rect -736 684 -731 687
rect -736 680 -711 684
rect -704 683 -700 697
rect -678 687 -671 730
rect -511 723 -470 731
rect -681 683 -671 687
rect -736 679 -728 680
rect -704 679 -677 683
rect -650 681 -646 700
rect -736 633 -731 679
rect -704 677 -700 679
rect -667 675 -646 681
rect -650 668 -646 675
rect -712 662 -708 667
rect -723 655 -687 662
rect -642 682 -638 700
rect -493 699 -488 711
rect -347 700 -343 705
rect -332 700 -328 769
rect -325 748 -322 752
rect -315 745 -311 776
rect -287 769 -283 776
rect -260 769 -256 776
rect -235 774 -231 825
rect -228 779 -224 838
rect -219 836 -191 839
rect -212 830 -209 836
rect -228 775 -211 779
rect -203 778 -200 790
rect -188 785 -147 788
rect -188 778 -185 785
rect -182 778 -154 781
rect -203 775 -185 778
rect -294 765 -283 769
rect -277 765 -256 769
rect -243 772 -231 774
rect -199 772 -195 775
rect -243 770 -195 772
rect -304 748 -301 752
rect -294 745 -290 765
rect -287 748 -284 752
rect -277 745 -273 765
rect -243 753 -239 770
rect -235 768 -195 770
rect -175 772 -172 778
rect -235 757 -207 760
rect -269 749 -266 753
rect -259 749 -239 753
rect -259 746 -255 749
rect -243 721 -239 749
rect -228 751 -225 757
rect -219 721 -216 731
rect -204 748 -174 751
rect -204 721 -201 748
rect -182 747 -174 748
rect -166 750 -163 762
rect -150 750 -147 785
rect -166 747 -147 750
rect -243 717 -227 721
rect -219 718 -201 721
rect -219 713 -216 718
rect -323 700 -319 705
rect -302 700 -298 705
rect -285 700 -281 705
rect -267 700 -263 706
rect -347 697 -263 700
rect -228 695 -225 703
rect -239 692 -225 695
rect -642 676 -607 682
rect -642 668 -638 676
rect -675 646 -649 653
rect -675 633 -668 646
rect -736 627 -668 633
rect -664 637 -656 641
rect -664 623 -661 637
rect -613 633 -607 676
rect -253 668 -225 671
rect -246 662 -243 668
rect -667 619 -661 623
rect -651 627 -607 633
rect -237 632 -234 642
rect -253 628 -245 632
rect -237 629 -225 632
rect -667 615 -664 619
rect -651 616 -647 627
rect -237 624 -234 629
rect -748 611 -664 615
rect -659 593 -655 606
rect -505 603 -498 612
rect -471 594 -464 610
rect -246 606 -243 614
rect -253 603 -243 606
rect 15 611 22 620
rect 49 602 56 618
rect -231 600 -228 602
rect -671 588 -635 593
rect -563 590 -464 594
rect -563 532 -554 590
rect -548 580 -505 587
rect -471 580 -464 590
rect -322 588 -319 592
rect -302 588 -296 592
rect -289 588 -286 592
rect -262 588 -259 592
rect -537 565 -533 580
rect -477 576 -450 580
rect -454 573 -450 576
rect -563 528 -536 532
rect -529 531 -525 545
rect -488 534 -484 553
rect -529 527 -502 531
rect -529 525 -525 527
rect -537 510 -533 515
rect -548 503 -512 510
rect -736 486 -662 491
rect -736 359 -730 486
rect -711 476 -678 483
rect -666 481 -662 486
rect -507 489 -502 527
rect -488 522 -484 528
rect -488 506 -484 512
rect -480 522 -476 553
rect -446 534 -442 553
rect -320 535 -316 544
rect -305 543 -300 544
rect -287 543 -283 545
rect -305 538 -283 543
rect -279 543 -275 545
rect -260 543 -256 545
rect -279 538 -256 543
rect -252 543 -248 545
rect -252 538 -243 543
rect -460 529 -453 533
rect -446 528 -423 534
rect -325 531 -307 535
rect -446 522 -442 528
rect -459 516 -454 522
rect -480 505 -476 512
rect -446 505 -442 512
rect -336 510 -333 514
rect -326 507 -322 516
rect -480 501 -442 505
rect -476 493 -472 498
rect -507 481 -466 489
rect -700 461 -696 476
rect -666 474 -637 481
rect -724 428 -719 431
rect -724 424 -699 428
rect -692 427 -688 441
rect -666 431 -659 474
rect -669 427 -659 431
rect -724 423 -716 424
rect -692 423 -665 427
rect -638 425 -634 444
rect -724 377 -719 423
rect -692 421 -688 423
rect -655 419 -634 425
rect -638 412 -634 419
rect -700 406 -696 411
rect -711 399 -675 406
rect -489 457 -484 469
rect -334 462 -330 467
rect -319 462 -315 531
rect -312 510 -309 514
rect -302 507 -298 538
rect -274 531 -270 538
rect -247 534 -243 538
rect -232 541 -228 600
rect -223 598 -195 601
rect -43 598 56 602
rect -216 592 -213 598
rect -232 537 -215 541
rect -207 540 -204 552
rect -192 547 -151 550
rect -192 540 -189 547
rect -186 540 -158 543
rect -207 537 -189 540
rect -203 534 -199 537
rect -281 527 -270 531
rect -264 530 -199 534
rect -179 534 -176 540
rect -291 510 -288 514
rect -281 507 -277 527
rect -274 510 -271 514
rect -264 507 -260 530
rect -247 483 -243 530
rect -239 519 -211 522
rect -232 513 -229 519
rect -223 483 -220 493
rect -208 510 -178 513
rect -208 483 -205 510
rect -186 509 -178 510
rect -170 512 -167 524
rect -154 512 -151 547
rect -43 540 -34 598
rect -28 588 15 595
rect 49 588 56 598
rect -17 573 -13 588
rect 43 584 70 588
rect 66 581 70 584
rect -43 536 -16 540
rect -9 539 -5 553
rect 32 542 36 561
rect -9 535 18 539
rect -9 533 -5 535
rect -17 518 -13 523
rect -170 509 -151 512
rect -28 511 8 518
rect 13 497 18 535
rect 32 530 36 536
rect 32 514 36 520
rect 40 530 44 561
rect 74 542 78 561
rect 60 537 67 541
rect 74 536 97 542
rect 74 530 78 536
rect 61 524 66 530
rect 40 513 44 520
rect 74 513 78 520
rect 40 509 78 513
rect 44 501 48 506
rect 13 489 54 497
rect -247 479 -231 483
rect -223 480 -205 483
rect -223 475 -220 480
rect -310 462 -306 467
rect -289 462 -285 467
rect -272 462 -268 467
rect 31 465 36 477
rect -334 459 -267 462
rect -232 457 -229 465
rect -243 454 -229 457
rect -630 426 -626 444
rect -248 441 -220 444
rect -241 435 -238 441
rect -630 420 -595 426
rect -630 412 -626 420
rect -663 390 -637 397
rect -663 377 -656 390
rect -724 371 -656 377
rect -652 381 -644 385
rect -652 367 -649 381
rect -601 377 -595 420
rect -232 405 -229 415
rect -248 401 -240 405
rect -232 402 -220 405
rect -232 397 -229 402
rect 19 389 26 398
rect -241 379 -238 387
rect 53 380 60 396
rect -655 363 -649 367
rect -639 371 -595 377
rect -655 359 -652 363
rect -639 360 -635 371
rect -493 369 -486 378
rect -248 376 -238 379
rect -39 376 60 380
rect -459 360 -452 376
rect -226 373 -223 375
rect -290 361 -287 365
rect -270 361 -264 365
rect -257 361 -254 365
rect -736 355 -652 359
rect -551 356 -452 360
rect -647 337 -643 350
rect -659 332 -623 337
rect -551 298 -542 356
rect -536 346 -493 353
rect -459 346 -452 356
rect -525 331 -521 346
rect -465 342 -438 346
rect -442 339 -438 342
rect -551 294 -524 298
rect -517 297 -513 311
rect -476 300 -472 319
rect -517 293 -490 297
rect -517 291 -513 293
rect -525 276 -521 281
rect -536 269 -500 276
rect -495 255 -490 293
rect -476 288 -472 294
rect -476 272 -472 278
rect -468 288 -464 319
rect -434 300 -430 319
rect -288 308 -284 317
rect -273 316 -268 317
rect -255 316 -251 318
rect -273 311 -251 316
rect -247 316 -243 318
rect -247 314 -241 316
rect -227 314 -223 373
rect -218 371 -190 374
rect -211 365 -208 371
rect -247 311 -239 314
rect -293 304 -275 308
rect -448 295 -441 299
rect -434 294 -411 300
rect -434 288 -430 294
rect -447 282 -442 288
rect -304 283 -301 287
rect -294 280 -290 289
rect -468 271 -464 278
rect -434 271 -430 278
rect -468 267 -430 271
rect -464 259 -460 264
rect -495 247 -454 255
rect -477 223 -472 235
rect -302 235 -298 240
rect -287 235 -283 304
rect -280 283 -277 287
rect -270 280 -266 311
rect -243 307 -239 311
rect -227 310 -210 314
rect -202 313 -199 325
rect -187 320 -146 323
rect -187 313 -184 320
rect -181 313 -153 316
rect -202 310 -184 313
rect -198 307 -194 310
rect -243 304 -194 307
rect -249 303 -194 304
rect -174 307 -171 313
rect -249 300 -236 303
rect -259 283 -256 287
rect -249 280 -245 300
rect -242 256 -238 300
rect -234 292 -206 295
rect -227 286 -224 292
rect -218 256 -215 266
rect -203 283 -173 286
rect -203 256 -200 283
rect -181 282 -173 283
rect -165 285 -162 297
rect -149 285 -146 320
rect -39 318 -30 376
rect -24 366 19 373
rect 53 366 60 376
rect -13 351 -9 366
rect 47 362 74 366
rect 70 359 74 362
rect -39 314 -12 318
rect -5 317 -1 331
rect 36 320 40 339
rect -5 313 22 317
rect -5 311 -1 313
rect -13 296 -9 301
rect -24 289 12 296
rect -165 282 -146 285
rect 17 275 22 313
rect 36 308 40 314
rect 36 292 40 298
rect 44 308 48 339
rect 78 320 82 339
rect 64 315 71 319
rect 78 314 101 320
rect 78 308 82 314
rect 65 302 70 308
rect 44 291 48 298
rect 78 291 82 298
rect 44 287 82 291
rect 48 279 52 284
rect 17 267 58 275
rect -242 252 -226 256
rect -218 253 -200 256
rect -218 248 -215 253
rect -278 235 -274 240
rect -257 235 -253 240
rect 35 243 40 255
rect -302 232 -243 235
rect -227 230 -224 238
rect -238 227 -224 230
rect -246 218 -218 221
rect -239 212 -236 218
rect -230 182 -227 192
rect -246 178 -238 182
rect -230 179 -218 182
rect -230 174 -227 179
rect 26 176 33 185
rect 60 167 67 183
rect -486 153 -479 162
rect -452 144 -445 160
rect -239 156 -236 164
rect -246 153 -236 156
rect -32 163 67 167
rect -224 150 -221 152
rect -544 140 -445 144
rect -713 111 -639 116
rect -713 -16 -707 111
rect -688 101 -655 108
rect -643 106 -639 111
rect -677 86 -673 101
rect -643 99 -614 106
rect -701 53 -696 56
rect -701 49 -676 53
rect -669 52 -665 66
rect -643 56 -636 99
rect -646 52 -636 56
rect -701 48 -693 49
rect -669 48 -642 52
rect -615 50 -611 69
rect -701 2 -696 48
rect -669 46 -665 48
rect -632 44 -611 50
rect -615 37 -611 44
rect -677 31 -673 36
rect -688 24 -652 31
rect -544 82 -535 140
rect -529 130 -486 137
rect -452 130 -445 140
rect -269 138 -266 142
rect -249 138 -243 142
rect -518 115 -514 130
rect -458 126 -431 130
rect -435 123 -431 126
rect -544 78 -517 82
rect -510 81 -506 95
rect -469 84 -465 103
rect -510 77 -483 81
rect -510 75 -506 77
rect -607 51 -603 69
rect -518 60 -514 65
rect -529 53 -493 60
rect -607 45 -572 51
rect -607 37 -603 45
rect -640 15 -614 22
rect -640 2 -633 15
rect -701 -4 -633 2
rect -629 6 -621 10
rect -629 -8 -626 6
rect -578 2 -572 45
rect -488 39 -483 77
rect -469 72 -465 78
rect -469 56 -465 62
rect -461 72 -457 103
rect -427 84 -423 103
rect -267 85 -263 94
rect -252 93 -247 94
rect -252 88 -246 93
rect -225 91 -221 150
rect -216 148 -188 151
rect -209 142 -206 148
rect -441 79 -434 83
rect -427 78 -404 84
rect -272 81 -254 85
rect -249 84 -245 88
rect -225 87 -208 91
rect -200 90 -197 102
rect -32 105 -23 163
rect -17 153 26 160
rect 60 153 67 163
rect -6 138 -2 153
rect 54 149 81 153
rect 77 146 81 149
rect -32 101 -5 105
rect 2 104 6 118
rect 43 107 47 126
rect 2 100 29 104
rect -185 97 -144 100
rect 2 98 6 100
rect -185 90 -182 97
rect -179 90 -151 93
rect -200 87 -182 90
rect -196 84 -192 87
rect -427 72 -423 78
rect -440 66 -435 72
rect -461 55 -457 62
rect -427 55 -423 62
rect -283 60 -280 64
rect -273 57 -269 66
rect -461 51 -423 55
rect -457 43 -453 48
rect -488 31 -447 39
rect -470 7 -465 19
rect -281 12 -277 17
rect -266 12 -262 81
rect -249 80 -192 84
rect -172 84 -169 90
rect -259 60 -256 64
rect -249 57 -245 80
rect -240 33 -236 80
rect -232 69 -204 72
rect -225 63 -222 69
rect -216 33 -213 43
rect -201 60 -171 63
rect -201 33 -198 60
rect -179 59 -171 60
rect -163 62 -160 74
rect -147 62 -144 97
rect -6 83 -2 88
rect -17 76 19 83
rect -163 59 -144 62
rect 24 62 29 100
rect 43 95 47 101
rect 43 79 47 85
rect 51 95 55 126
rect 85 107 89 126
rect 71 102 78 106
rect 85 101 108 107
rect 85 95 89 101
rect 72 89 77 95
rect 51 78 55 85
rect 85 78 89 85
rect 51 74 89 78
rect 55 66 59 71
rect 24 54 65 62
rect -240 29 -224 33
rect -216 30 -198 33
rect 42 30 47 42
rect -216 25 -213 30
rect -257 12 -253 17
rect -281 9 -239 12
rect -225 7 -222 15
rect -236 4 -222 7
rect -632 -12 -626 -8
rect -616 -4 -572 2
rect 35 3 42 12
rect -632 -16 -629 -12
rect -616 -15 -612 -4
rect 69 -6 76 10
rect -713 -20 -629 -16
rect -23 -10 76 -6
rect -624 -38 -620 -25
rect -636 -43 -600 -38
rect -23 -68 -14 -10
rect -8 -20 35 -13
rect 69 -20 76 -10
rect 3 -35 7 -20
rect 63 -24 90 -20
rect 86 -27 90 -24
rect -23 -72 4 -68
rect 11 -69 15 -55
rect 52 -66 56 -47
rect 11 -73 38 -69
rect 11 -75 15 -73
rect 3 -90 7 -85
rect -8 -97 28 -90
rect 33 -111 38 -73
rect 52 -78 56 -72
rect 52 -94 56 -88
rect 60 -78 64 -47
rect 94 -66 98 -47
rect 80 -71 87 -67
rect 94 -72 117 -66
rect 94 -78 98 -72
rect 81 -84 86 -78
rect 60 -95 64 -88
rect 94 -95 98 -88
rect 60 -99 98 -95
rect 64 -107 68 -102
rect 33 -119 74 -111
rect 51 -143 56 -131
<< m2contact >>
rect -509 839 -502 845
rect -509 822 -502 829
rect -493 770 -487 776
rect -493 743 -488 748
rect -469 770 -464 776
rect -470 758 -463 764
rect -476 735 -471 740
rect -470 723 -463 731
rect -493 711 -488 717
rect -505 597 -498 603
rect 15 605 22 611
rect -505 580 -498 587
rect -489 528 -483 534
rect -489 501 -484 506
rect -465 528 -460 534
rect -466 516 -459 522
rect -472 493 -467 498
rect -466 481 -459 489
rect -489 469 -484 475
rect 15 588 22 595
rect 31 536 37 542
rect 31 509 36 514
rect 55 536 60 542
rect 54 524 61 530
rect 48 501 53 506
rect 54 489 61 497
rect 31 477 36 483
rect 19 383 26 389
rect -493 363 -486 369
rect -493 346 -486 353
rect -477 294 -471 300
rect -477 267 -472 272
rect -453 294 -448 300
rect -454 282 -447 288
rect -460 259 -455 264
rect -454 247 -447 255
rect -477 235 -472 241
rect 19 366 26 373
rect 35 314 41 320
rect 35 287 40 292
rect 59 314 64 320
rect 58 302 65 308
rect 52 279 57 284
rect 58 267 65 275
rect 35 255 40 261
rect 26 170 33 176
rect -486 147 -479 153
rect -486 130 -479 137
rect -470 78 -464 84
rect -470 51 -465 56
rect -446 78 -441 84
rect 26 153 33 160
rect 42 101 48 107
rect -447 66 -440 72
rect -453 43 -448 48
rect -447 31 -440 39
rect -470 19 -465 25
rect 42 74 47 79
rect 66 101 71 107
rect 65 89 72 95
rect 59 66 64 71
rect 65 54 72 62
rect 42 42 47 48
rect 35 -3 42 3
rect 35 -20 42 -13
rect 51 -72 57 -66
rect 51 -99 56 -94
rect 75 -72 80 -66
rect 74 -84 81 -78
rect 68 -107 73 -102
rect 74 -119 81 -111
rect 51 -131 56 -125
<< metal2 >>
rect -509 829 -502 839
rect -487 771 -469 775
rect -493 717 -488 743
rect -470 740 -463 758
rect -471 735 -463 740
rect -470 731 -463 735
rect -505 587 -498 597
rect 15 595 22 605
rect 37 537 55 541
rect -483 529 -465 533
rect -489 475 -484 501
rect -466 498 -459 516
rect -467 493 -459 498
rect -466 489 -459 493
rect 31 483 36 509
rect 54 506 61 524
rect 53 501 61 506
rect 54 497 61 501
rect 19 373 26 383
rect -493 353 -486 363
rect 41 315 59 319
rect -471 295 -453 299
rect -477 241 -472 267
rect -454 264 -447 282
rect -455 259 -447 264
rect -454 255 -447 259
rect 35 261 40 287
rect 58 284 65 302
rect 57 279 65 284
rect 58 275 65 279
rect 26 160 33 170
rect -486 137 -479 147
rect 48 102 66 106
rect -464 79 -446 83
rect -470 25 -465 51
rect -447 48 -440 66
rect -448 43 -440 48
rect -447 39 -440 43
rect 42 48 47 74
rect 65 71 72 89
rect 64 66 72 71
rect 65 62 72 66
rect 35 -13 42 -3
rect 57 -71 75 -67
rect 51 -125 56 -99
rect 74 -102 81 -84
rect 73 -107 81 -102
rect 74 -111 81 -107
<< labels >>
rlabel metal1 -251 827 -250 828 1 p3
rlabel metal1 -274 827 -273 828 1 p2
rlabel metal1 -301 827 -300 828 1 p1
rlabel metal1 -334 827 -333 828 1 cin
rlabel metal1 -268 750 -267 751 1 g3
rlabel metal1 -286 749 -285 750 1 g2
rlabel metal1 -303 749 -302 750 1 g1
rlabel metal1 -324 749 -323 750 1 g0
rlabel metal1 -235 693 -233 694 1 gnd
rlabel metal1 -227 758 -225 759 1 vdd
rlabel metal1 -313 827 -312 829 1 p0
rlabel metal1 -169 779 -162 780 1 vdd
rlabel metal1 -206 837 -199 838 1 vdd
rlabel metal1 -241 907 -239 908 1 vdd
rlabel metal1 -249 842 -247 843 1 gnd
rlabel metal1 -219 775 -213 779 1 clk
rlabel metal1 -204 718 -201 751 1 c3
rlabel metal1 -242 825 -231 829 1 c3bar
rlabel metal1 -349 748 -346 752 3 clk
rlabel metal1 -339 745 -335 754 1 gnd
rlabel metal1 -249 866 -241 870 1 clk_org
rlabel metal1 -233 867 -221 870 1 clk
rlabel metal1 -239 455 -237 456 1 gnd
rlabel metal1 -231 520 -229 521 1 vdd
rlabel metal1 -173 541 -166 542 1 vdd
rlabel metal1 -210 599 -203 600 1 vdd
rlabel metal1 -245 669 -243 670 1 vdd
rlabel metal1 -253 604 -251 605 1 gnd
rlabel metal1 -223 537 -217 541 1 clk
rlabel metal1 -253 628 -245 632 1 clk_org
rlabel metal1 -237 629 -225 632 1 clk
rlabel metal1 -261 589 -260 590 1 p2
rlabel metal1 -288 589 -287 590 1 p1
rlabel metal1 -321 589 -320 590 1 cin
rlabel metal1 -273 511 -272 512 1 g2
rlabel metal1 -290 511 -289 512 1 g1
rlabel metal1 -311 511 -310 512 1 g0
rlabel metal1 -300 589 -299 591 1 p0
rlabel metal1 -336 510 -333 514 3 clk
rlabel metal1 -326 507 -322 516 1 gnd
rlabel metal1 -234 228 -232 229 1 gnd
rlabel metal1 -226 293 -224 294 1 vdd
rlabel metal1 -168 314 -161 315 1 vdd
rlabel metal1 -205 372 -198 373 1 vdd
rlabel metal1 -240 442 -238 443 1 vdd
rlabel metal1 -248 377 -246 378 1 gnd
rlabel metal1 -218 310 -212 314 1 clk
rlabel metal1 -248 401 -240 405 1 clk_org
rlabel metal1 -232 402 -220 405 1 clk
rlabel metal1 -247 479 -243 543 1 c2bar
rlabel metal1 -208 480 -205 513 1 c2
rlabel metal1 -294 280 -290 289 1 gnd
rlabel metal1 -304 283 -301 287 3 clk
rlabel metal1 -268 362 -267 364 1 p0
rlabel metal1 -279 284 -278 285 1 g0
rlabel metal1 -258 284 -257 285 1 g1
rlabel metal1 -289 362 -288 363 1 cin
rlabel metal1 -256 362 -255 363 1 p1
rlabel metal1 -243 300 -236 307 1 c1bar
rlabel metal1 -203 253 -200 286 1 c1
rlabel metal1 -232 5 -230 6 1 gnd
rlabel metal1 -224 70 -222 71 1 vdd
rlabel metal1 -166 91 -159 92 1 vdd
rlabel metal1 -203 149 -196 150 1 vdd
rlabel metal1 -238 219 -236 220 1 vdd
rlabel metal1 -246 154 -244 155 1 gnd
rlabel metal1 -216 87 -210 91 1 clk
rlabel metal1 -246 178 -238 182 1 clk_org
rlabel metal1 -230 179 -218 182 1 clk
rlabel metal1 -273 57 -269 66 1 gnd
rlabel metal1 -283 60 -280 64 3 clk
rlabel metal1 -247 139 -246 141 1 p0
rlabel metal1 -258 61 -257 62 1 g0
rlabel metal1 -268 139 -267 140 1 cin
rlabel metal1 -249 80 -192 84 1 c0bar
rlabel metal1 -201 30 -198 63 1 c0
rlabel metal1 -8 592 -8 592 1 vdd
rlabel metal1 -7 512 -7 512 1 gnd
rlabel metal1 18 616 18 616 5 vdd
rlabel metal1 -8 514 -8 514 1 gnd
rlabel metal1 -9 592 -9 592 5 vdd
rlabel metal1 -4 370 -4 370 1 vdd
rlabel metal1 -3 290 -3 290 1 gnd
rlabel metal1 22 394 22 394 5 vdd
rlabel metal1 -4 292 -4 292 1 gnd
rlabel metal1 -5 370 -5 370 5 vdd
rlabel metal1 3 157 3 157 1 vdd
rlabel metal1 4 77 4 77 1 gnd
rlabel metal1 29 181 29 181 5 vdd
rlabel metal1 3 79 3 79 1 gnd
rlabel metal1 2 157 2 157 5 vdd
rlabel metal1 -532 826 -532 826 1 vdd
rlabel metal1 -531 746 -531 746 1 gnd
rlabel metal1 -506 850 -506 850 5 vdd
rlabel metal1 -532 748 -532 748 1 gnd
rlabel metal1 -533 826 -533 826 5 vdd
rlabel metal1 -528 584 -528 584 1 vdd
rlabel metal1 -527 504 -527 504 1 gnd
rlabel metal1 -502 608 -502 608 5 vdd
rlabel metal1 -528 506 -528 506 1 gnd
rlabel metal1 -529 584 -529 584 5 vdd
rlabel metal1 -516 350 -516 350 1 vdd
rlabel metal1 -515 270 -515 270 1 gnd
rlabel metal1 -490 374 -490 374 5 vdd
rlabel metal1 -516 272 -516 272 1 gnd
rlabel metal1 -517 350 -517 350 5 vdd
rlabel metal1 -510 134 -510 134 5 vdd
rlabel metal1 -509 56 -509 56 1 gnd
rlabel metal1 -483 158 -483 158 5 vdd
rlabel metal1 -508 54 -508 54 1 gnd
rlabel metal1 -509 134 -509 134 1 vdd
rlabel metal1 11 -16 11 -16 5 vdd
rlabel metal1 12 -94 12 -94 1 gnd
rlabel metal1 38 8 38 8 5 vdd
rlabel metal1 13 -96 13 -96 1 gnd
rlabel metal1 12 -16 12 -16 1 vdd
rlabel metal1 31 465 36 477 1 p3
rlabel metal1 49 584 56 618 1 c2
rlabel metal1 35 243 40 255 1 p2
rlabel metal1 53 362 60 396 1 c1
rlabel metal1 42 30 47 42 1 p1
rlabel metal1 -32 163 67 167 1 c0
rlabel metal1 51 -143 56 -131 1 p0
rlabel metal1 69 -24 76 10 1 cin
rlabel metal1 -470 7 -465 19 1 a0
rlabel metal1 -477 223 -472 235 1 a1
rlabel metal1 -459 342 -452 376 1 b1
rlabel metal1 -489 457 -484 469 1 a2
rlabel metal1 -471 576 -464 610 1 b2
rlabel metal1 -493 699 -488 711 1 a3
rlabel metal1 -475 818 -468 852 1 b3
rlabel metal1 -704 736 -704 736 5 vdd
rlabel metal1 -703 658 -703 658 1 gnd
rlabel metal1 -658 590 -658 590 1 gnd
rlabel metal1 -692 480 -692 480 5 vdd
rlabel metal1 -691 402 -691 402 1 gnd
rlabel metal1 -646 334 -646 334 1 gnd
rlabel metal1 -669 105 -669 105 5 vdd
rlabel metal1 -668 27 -668 27 1 gnd
rlabel metal1 -623 -41 -623 -41 1 gnd
rlabel metal1 -710 1020 -710 1020 5 vdd
rlabel metal1 -709 942 -709 942 1 gnd
rlabel metal1 -664 874 -664 874 1 gnd
rlabel metal1 -742 911 -737 971 1 a3
rlabel metal1 -673 959 -652 965 1 b3
rlabel metal1 -736 627 -731 687 1 a2
rlabel metal1 -667 675 -646 681 1 b2
rlabel metal1 -724 371 -719 431 1 a1
rlabel metal1 -655 419 -634 425 1 b1
rlabel metal1 -701 -4 -696 56 1 a0
rlabel metal1 -632 44 -611 50 1 b0
rlabel metal1 -619 911 -613 966 1 g3
rlabel metal1 -613 627 -607 682 1 g2
rlabel metal1 -601 371 -595 426 1 g1
rlabel metal1 -578 -4 -572 51 1 g0
rlabel metal1 -450 770 -427 776 1 p3
rlabel metal1 -446 528 -423 534 1 p2
rlabel metal1 -434 294 -411 300 1 p1
rlabel metal1 -427 78 -404 84 1 p0
rlabel metal1 74 536 97 542 1 s3in
rlabel metal1 78 314 101 320 1 s2in
rlabel metal1 85 101 108 107 1 s1in
rlabel metal1 94 -72 117 -66 1 s0in
<< end >>
