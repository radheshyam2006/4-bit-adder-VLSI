
.include TSMC_180nm.txt
.param SUPPLY=1.8
.param LAMBDA=0.09u

vdd vdd gnd DC 1.8

.subckt nmos d g s b W='N'
.param width_N={W}
M1 d g s b CMOSN W={width_N} L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N}
+ AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
.ends nmos

.subckt pmos d g s b W='P'
.param width_P={W}
M1 d g s b CMOSP W={width_P} L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P}
+ AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends pmos

.subckt inv out in vdd gnd N='a'
.param width_N={N}
.param width_P={2*width_N}
M1      out       in      gnd     gnd  CMOSN   W={width_N}   L={2*LAMBDA}
+ AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
M2      out       in      vdd     vdd  CMOSP   W={width_P}   L={2*LAMBDA}
+ AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends inv

* Logic gates and connections for the circuit
x1 n12 abar vdd vdd pmos W='20*LAMBDA'
x2 n23 bbar n12 n12 pmos W='20*LAMBDA'
x3 n67 a vdd vdd pmos W='20*LAMBDA'
x4 n23 b n67 n67 pmos W='20*LAMBDA'
x5 n34 clk n23 n23 pmos W='20*LAMBDA'
x6 n34 abar n45 n45 nmos W='10*LAMBDA'
x7 n45 b gnd gnd nmos W='10*LAMBDA'
x8 n34 a n89 n89 nmos W='10*LAMBDA'
x9 n89 bbar gnd gnd nmos W='10*LAMBDA'

x10 m67 n34 vdd vdd pmos W='20*LAMBDA'
x11 m78 clk m67 m67 pmos W='20*LAMBDA'
x12 m78 n34 gnd gnd nmos W='10*LAMBDA'

x13 m910 m78 vdd vdd pmos W='20*LAMBDA'
x14 m910 clk m1011 m1011 nmos W='10*LAMBDA'
x15 m1011 m78 gnd gnd nmos W='10*LAMBDA'

x16 out m910 vdd vdd pmos W='20*LAMBDA'
x17 out clk m1314 m1314 nmos W='10*LAMBDA'
x18 m1314 m910 gnd gnd nmos W='10*LAMBDA'

x19 abar a vdd gnd inv N='10*LAMBDA'
x20 bbar b vdd gnd inv N='10*LAMBDA'

* Stimuli
V1 clk gnd pulse(0 1.8 80n 0 0 40n 80n)
V2 a gnd pulse(0 1.8 10n 0 0 160n 320n)
V3 b gnd pulse(0 1.8 15n 0 0 320n 640n)

* Simulation settings
.tran 0.1n 640ns
.control
run
set hcopypscolor = 1
set color0 = white
set color1 = blue
plot v(clk) v(a)+6 v(b)+4 v(out)+2
.endc
