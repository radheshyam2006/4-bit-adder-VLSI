magic
tech scmos
timestamp 1732102597
<< nwell >>
rect 467 2215 504 2241
rect 510 2215 538 2241
rect 816 2236 850 2264
rect 458 2128 482 2152
rect 497 2142 531 2148
rect 497 2112 559 2142
rect 661 2136 689 2170
rect 819 2164 847 2218
rect 525 2106 559 2112
rect 803 2105 831 2139
rect 856 2136 884 2160
rect 458 2073 482 2097
rect 909 2042 933 2066
rect 948 2056 982 2062
rect 458 1980 495 2006
rect 501 1980 529 2006
rect 812 2002 846 2030
rect 948 2026 1010 2056
rect 976 2020 1010 2026
rect 456 1893 480 1917
rect 674 1913 702 1947
rect 815 1942 843 1996
rect 909 1987 933 2011
rect 495 1907 529 1913
rect 495 1877 557 1907
rect 799 1883 827 1917
rect 852 1914 880 1938
rect 523 1871 557 1877
rect 456 1838 480 1862
rect 908 1850 932 1874
rect 947 1864 981 1870
rect 817 1809 851 1837
rect 947 1834 1009 1864
rect 975 1828 1009 1834
rect 466 1761 503 1787
rect 509 1761 537 1787
rect 707 1719 735 1753
rect 820 1748 848 1802
rect 908 1795 932 1819
rect 453 1690 477 1714
rect 492 1704 526 1710
rect 492 1674 554 1704
rect 804 1689 832 1723
rect 857 1720 885 1744
rect 520 1668 554 1674
rect 453 1635 477 1659
rect 926 1653 950 1677
rect 965 1667 999 1673
rect 965 1637 1027 1667
rect 993 1631 1027 1637
rect 464 1569 501 1595
rect 507 1569 535 1595
rect 819 1571 853 1599
rect 926 1598 950 1622
rect 452 1494 476 1518
rect 491 1508 525 1514
rect 491 1478 553 1508
rect 726 1482 754 1516
rect 822 1510 850 1564
rect 519 1472 553 1478
rect 452 1439 476 1463
rect 806 1451 834 1485
rect 859 1482 887 1506
rect 687 1379 711 1403
rect 726 1393 760 1399
rect 726 1363 788 1393
rect 754 1357 788 1363
rect 687 1324 711 1348
<< ntransistor >>
rect 796 2250 806 2252
rect 480 2187 482 2200
rect 490 2187 492 2200
rect 522 2198 524 2205
rect 710 2164 712 2205
rect 717 2164 719 2205
rect 743 2165 745 2205
rect 770 2165 772 2205
rect 793 2165 795 2205
rect 469 2114 471 2120
rect 673 2116 675 2126
rect 696 2087 698 2127
rect 720 2087 722 2127
rect 741 2087 743 2127
rect 758 2087 760 2127
rect 776 2088 778 2128
rect 815 2085 817 2095
rect 508 2065 510 2077
rect 518 2065 520 2077
rect 536 2065 538 2077
rect 546 2065 548 2077
rect 469 2059 471 2065
rect 920 2028 922 2034
rect 792 2016 802 2018
rect 471 1952 473 1965
rect 481 1952 483 1965
rect 513 1963 515 1970
rect 723 1942 725 1983
rect 730 1942 732 1983
rect 756 1943 758 1983
rect 783 1943 785 1983
rect 959 1979 961 1991
rect 969 1979 971 1991
rect 987 1979 989 1991
rect 997 1979 999 1991
rect 920 1973 922 1979
rect 467 1879 469 1885
rect 686 1893 688 1903
rect 709 1865 711 1905
rect 733 1865 735 1905
rect 754 1865 756 1905
rect 771 1865 773 1905
rect 811 1863 813 1873
rect 506 1830 508 1842
rect 516 1830 518 1842
rect 534 1830 536 1842
rect 544 1830 546 1842
rect 919 1836 921 1842
rect 467 1824 469 1830
rect 797 1823 807 1825
rect 479 1733 481 1746
rect 489 1733 491 1746
rect 521 1744 523 1751
rect 755 1748 757 1789
rect 762 1748 764 1789
rect 788 1749 790 1789
rect 958 1787 960 1799
rect 968 1787 970 1799
rect 986 1787 988 1799
rect 996 1787 998 1799
rect 919 1781 921 1787
rect 464 1676 466 1682
rect 719 1699 721 1709
rect 741 1671 743 1711
rect 765 1671 767 1711
rect 786 1671 788 1711
rect 816 1669 818 1679
rect 937 1639 939 1645
rect 503 1627 505 1639
rect 513 1627 515 1639
rect 531 1627 533 1639
rect 541 1627 543 1639
rect 464 1621 466 1627
rect 976 1590 978 1602
rect 986 1590 988 1602
rect 1004 1590 1006 1602
rect 1014 1590 1016 1602
rect 799 1585 809 1587
rect 937 1584 939 1590
rect 477 1541 479 1554
rect 487 1541 489 1554
rect 519 1552 521 1559
rect 776 1510 778 1551
rect 783 1510 785 1551
rect 463 1480 465 1486
rect 738 1462 740 1472
rect 502 1431 504 1443
rect 512 1431 514 1443
rect 530 1431 532 1443
rect 540 1431 542 1443
rect 762 1433 764 1473
rect 786 1433 788 1473
rect 463 1425 465 1431
rect 818 1431 820 1441
rect 698 1365 700 1371
rect 737 1316 739 1328
rect 747 1316 749 1328
rect 765 1316 767 1328
rect 775 1316 777 1328
rect 698 1310 700 1316
<< ptransistor >>
rect 824 2250 844 2252
rect 480 2223 482 2235
rect 490 2223 492 2235
rect 522 2223 524 2235
rect 831 2172 833 2212
rect 469 2134 471 2146
rect 673 2144 675 2164
rect 868 2144 870 2154
rect 508 2118 510 2142
rect 518 2118 520 2142
rect 536 2112 538 2136
rect 546 2112 548 2136
rect 469 2079 471 2091
rect 815 2113 817 2133
rect 920 2048 922 2060
rect 959 2032 961 2056
rect 969 2032 971 2056
rect 987 2026 989 2050
rect 997 2026 999 2050
rect 820 2016 840 2018
rect 471 1988 473 2000
rect 481 1988 483 2000
rect 513 1988 515 2000
rect 920 1993 922 2005
rect 827 1950 829 1990
rect 686 1921 688 1941
rect 864 1922 866 1932
rect 467 1899 469 1911
rect 506 1883 508 1907
rect 516 1883 518 1907
rect 534 1877 536 1901
rect 544 1877 546 1901
rect 467 1844 469 1856
rect 811 1891 813 1911
rect 919 1856 921 1868
rect 958 1840 960 1864
rect 968 1840 970 1864
rect 986 1834 988 1858
rect 996 1834 998 1858
rect 825 1823 845 1825
rect 919 1801 921 1813
rect 479 1769 481 1781
rect 489 1769 491 1781
rect 521 1769 523 1781
rect 832 1756 834 1796
rect 719 1727 721 1747
rect 869 1728 871 1738
rect 464 1696 466 1708
rect 503 1680 505 1704
rect 513 1680 515 1704
rect 531 1674 533 1698
rect 541 1674 543 1698
rect 464 1641 466 1653
rect 816 1697 818 1717
rect 937 1659 939 1671
rect 976 1643 978 1667
rect 986 1643 988 1667
rect 1004 1637 1006 1661
rect 1014 1637 1016 1661
rect 937 1604 939 1616
rect 477 1577 479 1589
rect 487 1577 489 1589
rect 519 1577 521 1589
rect 827 1585 847 1587
rect 463 1500 465 1512
rect 834 1518 836 1558
rect 502 1484 504 1508
rect 512 1484 514 1508
rect 530 1478 532 1502
rect 540 1478 542 1502
rect 738 1490 740 1510
rect 871 1490 873 1500
rect 463 1445 465 1457
rect 818 1459 820 1479
rect 698 1385 700 1397
rect 737 1369 739 1393
rect 747 1369 749 1393
rect 765 1363 767 1387
rect 775 1363 777 1387
rect 698 1330 700 1342
<< ndiffusion >>
rect 796 2252 806 2253
rect 796 2249 806 2250
rect 479 2187 480 2200
rect 482 2187 490 2200
rect 492 2187 493 2200
rect 521 2198 522 2205
rect 524 2198 525 2205
rect 709 2164 710 2205
rect 712 2164 717 2205
rect 719 2164 720 2205
rect 742 2165 743 2205
rect 745 2165 746 2205
rect 769 2165 770 2205
rect 772 2165 773 2205
rect 792 2165 793 2205
rect 795 2165 796 2205
rect 468 2114 469 2120
rect 471 2114 472 2120
rect 672 2116 673 2126
rect 675 2116 676 2126
rect 695 2087 696 2127
rect 698 2087 699 2127
rect 719 2087 720 2127
rect 722 2087 723 2127
rect 740 2087 741 2127
rect 743 2087 744 2127
rect 757 2087 758 2127
rect 760 2087 761 2127
rect 775 2088 776 2128
rect 778 2088 779 2128
rect 814 2085 815 2095
rect 817 2085 818 2095
rect 507 2065 508 2077
rect 510 2065 518 2077
rect 520 2065 521 2077
rect 535 2065 536 2077
rect 538 2065 546 2077
rect 548 2065 549 2077
rect 468 2059 469 2065
rect 471 2059 472 2065
rect 919 2028 920 2034
rect 922 2028 923 2034
rect 792 2018 802 2019
rect 792 2015 802 2016
rect 470 1952 471 1965
rect 473 1952 481 1965
rect 483 1952 484 1965
rect 512 1963 513 1970
rect 515 1963 516 1970
rect 722 1942 723 1983
rect 725 1942 730 1983
rect 732 1942 733 1983
rect 755 1943 756 1983
rect 758 1943 759 1983
rect 782 1943 783 1983
rect 785 1943 786 1983
rect 958 1979 959 1991
rect 961 1979 969 1991
rect 971 1979 972 1991
rect 986 1979 987 1991
rect 989 1979 997 1991
rect 999 1979 1000 1991
rect 919 1973 920 1979
rect 922 1973 923 1979
rect 466 1879 467 1885
rect 469 1879 470 1885
rect 685 1893 686 1903
rect 688 1893 689 1903
rect 708 1865 709 1905
rect 711 1865 712 1905
rect 732 1865 733 1905
rect 735 1865 736 1905
rect 753 1865 754 1905
rect 756 1865 757 1905
rect 770 1865 771 1905
rect 773 1865 774 1905
rect 810 1863 811 1873
rect 813 1863 814 1873
rect 505 1830 506 1842
rect 508 1830 516 1842
rect 518 1830 519 1842
rect 533 1830 534 1842
rect 536 1830 544 1842
rect 546 1830 547 1842
rect 918 1836 919 1842
rect 921 1836 922 1842
rect 466 1824 467 1830
rect 469 1824 470 1830
rect 797 1825 807 1826
rect 797 1822 807 1823
rect 478 1733 479 1746
rect 481 1733 489 1746
rect 491 1733 492 1746
rect 520 1744 521 1751
rect 523 1744 524 1751
rect 754 1748 755 1789
rect 757 1748 762 1789
rect 764 1748 765 1789
rect 787 1749 788 1789
rect 790 1749 791 1789
rect 957 1787 958 1799
rect 960 1787 968 1799
rect 970 1787 971 1799
rect 985 1787 986 1799
rect 988 1787 996 1799
rect 998 1787 999 1799
rect 918 1781 919 1787
rect 921 1781 922 1787
rect 463 1676 464 1682
rect 466 1676 467 1682
rect 718 1699 719 1709
rect 721 1699 722 1709
rect 740 1671 741 1711
rect 743 1671 744 1711
rect 764 1671 765 1711
rect 767 1671 768 1711
rect 785 1671 786 1711
rect 788 1671 789 1711
rect 815 1669 816 1679
rect 818 1669 819 1679
rect 936 1639 937 1645
rect 939 1639 940 1645
rect 502 1627 503 1639
rect 505 1627 513 1639
rect 515 1627 516 1639
rect 530 1627 531 1639
rect 533 1627 541 1639
rect 543 1627 544 1639
rect 463 1621 464 1627
rect 466 1621 467 1627
rect 799 1587 809 1588
rect 975 1590 976 1602
rect 978 1590 986 1602
rect 988 1590 989 1602
rect 1003 1590 1004 1602
rect 1006 1590 1014 1602
rect 1016 1590 1017 1602
rect 799 1584 809 1585
rect 936 1584 937 1590
rect 939 1584 940 1590
rect 476 1541 477 1554
rect 479 1541 487 1554
rect 489 1541 490 1554
rect 518 1552 519 1559
rect 521 1552 522 1559
rect 775 1510 776 1551
rect 778 1510 783 1551
rect 785 1510 786 1551
rect 462 1480 463 1486
rect 465 1480 466 1486
rect 737 1462 738 1472
rect 740 1462 741 1472
rect 501 1431 502 1443
rect 504 1431 512 1443
rect 514 1431 515 1443
rect 529 1431 530 1443
rect 532 1431 540 1443
rect 542 1431 543 1443
rect 761 1433 762 1473
rect 764 1433 765 1473
rect 785 1433 786 1473
rect 788 1433 789 1473
rect 462 1425 463 1431
rect 465 1425 466 1431
rect 817 1431 818 1441
rect 820 1431 821 1441
rect 697 1365 698 1371
rect 700 1365 701 1371
rect 736 1316 737 1328
rect 739 1316 747 1328
rect 749 1316 750 1328
rect 764 1316 765 1328
rect 767 1316 775 1328
rect 777 1316 778 1328
rect 697 1310 698 1316
rect 700 1310 701 1316
<< pdiffusion >>
rect 824 2252 844 2253
rect 824 2249 844 2250
rect 479 2223 480 2235
rect 482 2223 484 2235
rect 488 2223 490 2235
rect 492 2223 493 2235
rect 521 2223 522 2235
rect 524 2223 525 2235
rect 830 2172 831 2212
rect 833 2172 834 2212
rect 468 2134 469 2146
rect 471 2134 472 2146
rect 672 2144 673 2164
rect 675 2144 676 2164
rect 867 2144 868 2154
rect 870 2144 871 2154
rect 507 2118 508 2142
rect 510 2118 512 2142
rect 516 2118 518 2142
rect 520 2118 521 2142
rect 535 2112 536 2136
rect 538 2112 540 2136
rect 544 2112 546 2136
rect 548 2112 549 2136
rect 468 2079 469 2091
rect 471 2079 472 2091
rect 814 2113 815 2133
rect 817 2113 818 2133
rect 919 2048 920 2060
rect 922 2048 923 2060
rect 958 2032 959 2056
rect 961 2032 963 2056
rect 967 2032 969 2056
rect 971 2032 972 2056
rect 820 2018 840 2019
rect 986 2026 987 2050
rect 989 2026 991 2050
rect 995 2026 997 2050
rect 999 2026 1000 2050
rect 820 2015 840 2016
rect 470 1988 471 2000
rect 473 1988 475 2000
rect 479 1988 481 2000
rect 483 1988 484 2000
rect 512 1988 513 2000
rect 515 1988 516 2000
rect 919 1993 920 2005
rect 922 1993 923 2005
rect 826 1950 827 1990
rect 829 1950 830 1990
rect 685 1921 686 1941
rect 688 1921 689 1941
rect 863 1922 864 1932
rect 866 1922 867 1932
rect 466 1899 467 1911
rect 469 1899 470 1911
rect 505 1883 506 1907
rect 508 1883 510 1907
rect 514 1883 516 1907
rect 518 1883 519 1907
rect 533 1877 534 1901
rect 536 1877 538 1901
rect 542 1877 544 1901
rect 546 1877 547 1901
rect 466 1844 467 1856
rect 469 1844 470 1856
rect 810 1891 811 1911
rect 813 1891 814 1911
rect 918 1856 919 1868
rect 921 1856 922 1868
rect 957 1840 958 1864
rect 960 1840 962 1864
rect 966 1840 968 1864
rect 970 1840 971 1864
rect 985 1834 986 1858
rect 988 1834 990 1858
rect 994 1834 996 1858
rect 998 1834 999 1858
rect 825 1825 845 1826
rect 825 1822 845 1823
rect 918 1801 919 1813
rect 921 1801 922 1813
rect 478 1769 479 1781
rect 481 1769 483 1781
rect 487 1769 489 1781
rect 491 1769 492 1781
rect 520 1769 521 1781
rect 523 1769 524 1781
rect 831 1756 832 1796
rect 834 1756 835 1796
rect 718 1727 719 1747
rect 721 1727 722 1747
rect 868 1728 869 1738
rect 871 1728 872 1738
rect 463 1696 464 1708
rect 466 1696 467 1708
rect 502 1680 503 1704
rect 505 1680 507 1704
rect 511 1680 513 1704
rect 515 1680 516 1704
rect 530 1674 531 1698
rect 533 1674 535 1698
rect 539 1674 541 1698
rect 543 1674 544 1698
rect 463 1641 464 1653
rect 466 1641 467 1653
rect 815 1697 816 1717
rect 818 1697 819 1717
rect 936 1659 937 1671
rect 939 1659 940 1671
rect 975 1643 976 1667
rect 978 1643 980 1667
rect 984 1643 986 1667
rect 988 1643 989 1667
rect 1003 1637 1004 1661
rect 1006 1637 1008 1661
rect 1012 1637 1014 1661
rect 1016 1637 1017 1661
rect 936 1604 937 1616
rect 939 1604 940 1616
rect 476 1577 477 1589
rect 479 1577 481 1589
rect 485 1577 487 1589
rect 489 1577 490 1589
rect 518 1577 519 1589
rect 521 1577 522 1589
rect 827 1587 847 1588
rect 827 1584 847 1585
rect 462 1500 463 1512
rect 465 1500 466 1512
rect 833 1518 834 1558
rect 836 1518 837 1558
rect 501 1484 502 1508
rect 504 1484 506 1508
rect 510 1484 512 1508
rect 514 1484 515 1508
rect 529 1478 530 1502
rect 532 1478 534 1502
rect 538 1478 540 1502
rect 542 1478 543 1502
rect 737 1490 738 1510
rect 740 1490 741 1510
rect 870 1490 871 1500
rect 873 1490 874 1500
rect 462 1445 463 1457
rect 465 1445 466 1457
rect 817 1459 818 1479
rect 820 1459 821 1479
rect 697 1385 698 1397
rect 700 1385 701 1397
rect 736 1369 737 1393
rect 739 1369 741 1393
rect 745 1369 747 1393
rect 749 1369 750 1393
rect 764 1363 765 1387
rect 767 1363 769 1387
rect 773 1363 775 1387
rect 777 1363 778 1387
rect 697 1330 698 1342
rect 700 1330 701 1342
<< ndcontact >>
rect 796 2253 806 2257
rect 796 2245 806 2249
rect 475 2187 479 2200
rect 493 2187 497 2200
rect 517 2198 521 2205
rect 525 2198 529 2205
rect 705 2164 709 2205
rect 720 2164 725 2205
rect 738 2165 742 2205
rect 746 2165 750 2205
rect 765 2165 769 2205
rect 773 2165 777 2205
rect 788 2165 792 2205
rect 796 2165 800 2205
rect 464 2114 468 2120
rect 472 2114 476 2120
rect 668 2116 672 2126
rect 676 2116 680 2126
rect 691 2087 695 2127
rect 699 2087 703 2127
rect 715 2087 719 2127
rect 723 2087 727 2127
rect 736 2087 740 2127
rect 744 2087 748 2127
rect 753 2087 757 2127
rect 761 2087 765 2127
rect 771 2088 775 2128
rect 779 2088 783 2128
rect 810 2085 814 2095
rect 818 2085 822 2095
rect 503 2065 507 2077
rect 521 2065 525 2077
rect 531 2065 535 2077
rect 549 2065 553 2077
rect 464 2059 468 2065
rect 472 2059 476 2065
rect 915 2028 919 2034
rect 923 2028 927 2034
rect 792 2019 802 2023
rect 792 2011 802 2015
rect 466 1952 470 1965
rect 484 1952 488 1965
rect 508 1963 512 1970
rect 516 1963 520 1970
rect 718 1942 722 1983
rect 733 1942 738 1983
rect 751 1943 755 1983
rect 759 1943 763 1983
rect 778 1943 782 1983
rect 786 1943 790 1983
rect 954 1979 958 1991
rect 972 1979 976 1991
rect 982 1979 986 1991
rect 1000 1979 1004 1991
rect 915 1973 919 1979
rect 923 1973 927 1979
rect 462 1879 466 1885
rect 470 1879 474 1885
rect 681 1893 685 1903
rect 689 1893 693 1903
rect 704 1865 708 1905
rect 712 1865 716 1905
rect 728 1865 732 1905
rect 736 1865 740 1905
rect 749 1865 753 1905
rect 757 1865 761 1905
rect 766 1865 770 1905
rect 774 1865 778 1905
rect 806 1863 810 1873
rect 814 1863 818 1873
rect 501 1830 505 1842
rect 519 1830 523 1842
rect 529 1830 533 1842
rect 547 1830 551 1842
rect 914 1836 918 1842
rect 922 1836 926 1842
rect 462 1824 466 1830
rect 470 1824 474 1830
rect 797 1826 807 1830
rect 797 1818 807 1822
rect 474 1733 478 1746
rect 492 1733 496 1746
rect 516 1744 520 1751
rect 524 1744 528 1751
rect 750 1748 754 1789
rect 765 1748 770 1789
rect 783 1749 787 1789
rect 791 1749 795 1789
rect 953 1787 957 1799
rect 971 1787 975 1799
rect 981 1787 985 1799
rect 999 1787 1003 1799
rect 914 1781 918 1787
rect 922 1781 926 1787
rect 459 1676 463 1682
rect 467 1676 471 1682
rect 714 1699 718 1709
rect 722 1699 726 1709
rect 736 1671 740 1711
rect 744 1671 748 1711
rect 760 1671 764 1711
rect 768 1671 772 1711
rect 781 1671 785 1711
rect 789 1671 793 1711
rect 811 1669 815 1679
rect 819 1669 823 1679
rect 932 1639 936 1645
rect 940 1639 944 1645
rect 498 1627 502 1639
rect 516 1627 520 1639
rect 526 1627 530 1639
rect 544 1627 548 1639
rect 459 1621 463 1627
rect 467 1621 471 1627
rect 799 1588 809 1592
rect 971 1590 975 1602
rect 989 1590 993 1602
rect 999 1590 1003 1602
rect 1017 1590 1021 1602
rect 799 1580 809 1584
rect 932 1584 936 1590
rect 940 1584 944 1590
rect 472 1541 476 1554
rect 490 1541 494 1554
rect 514 1552 518 1559
rect 522 1552 526 1559
rect 771 1510 775 1551
rect 786 1510 791 1551
rect 458 1480 462 1486
rect 466 1480 470 1486
rect 733 1462 737 1472
rect 741 1462 745 1472
rect 497 1431 501 1443
rect 515 1431 519 1443
rect 525 1431 529 1443
rect 543 1431 547 1443
rect 757 1433 761 1473
rect 765 1433 769 1473
rect 781 1433 785 1473
rect 789 1433 793 1473
rect 458 1425 462 1431
rect 466 1425 470 1431
rect 813 1431 817 1441
rect 821 1431 825 1441
rect 693 1365 697 1371
rect 701 1365 705 1371
rect 732 1316 736 1328
rect 750 1316 754 1328
rect 760 1316 764 1328
rect 778 1316 782 1328
rect 693 1310 697 1316
rect 701 1310 705 1316
<< pdcontact >>
rect 824 2253 844 2257
rect 824 2245 844 2249
rect 475 2223 479 2235
rect 484 2223 488 2235
rect 493 2223 497 2235
rect 517 2223 521 2235
rect 525 2223 529 2235
rect 826 2172 830 2212
rect 834 2172 838 2212
rect 464 2134 468 2146
rect 472 2134 476 2146
rect 668 2144 672 2164
rect 676 2144 680 2164
rect 863 2144 867 2154
rect 871 2144 875 2154
rect 503 2118 507 2142
rect 512 2118 516 2142
rect 521 2118 525 2142
rect 531 2112 535 2136
rect 540 2112 544 2136
rect 549 2112 553 2136
rect 464 2079 468 2091
rect 472 2079 476 2091
rect 810 2113 814 2133
rect 818 2113 822 2133
rect 915 2048 919 2060
rect 923 2048 927 2060
rect 954 2032 958 2056
rect 963 2032 967 2056
rect 972 2032 976 2056
rect 820 2019 840 2023
rect 982 2026 986 2050
rect 991 2026 995 2050
rect 1000 2026 1004 2050
rect 820 2011 840 2015
rect 466 1988 470 2000
rect 475 1988 479 2000
rect 484 1988 488 2000
rect 508 1988 512 2000
rect 516 1988 520 2000
rect 915 1993 919 2005
rect 923 1993 927 2005
rect 822 1950 826 1990
rect 830 1950 834 1990
rect 681 1921 685 1941
rect 689 1921 693 1941
rect 859 1922 863 1932
rect 867 1922 871 1932
rect 462 1899 466 1911
rect 470 1899 474 1911
rect 501 1883 505 1907
rect 510 1883 514 1907
rect 519 1883 523 1907
rect 529 1877 533 1901
rect 538 1877 542 1901
rect 547 1877 551 1901
rect 462 1844 466 1856
rect 470 1844 474 1856
rect 806 1891 810 1911
rect 814 1891 818 1911
rect 914 1856 918 1868
rect 922 1856 926 1868
rect 953 1840 957 1864
rect 962 1840 966 1864
rect 971 1840 975 1864
rect 825 1826 845 1830
rect 981 1834 985 1858
rect 990 1834 994 1858
rect 999 1834 1003 1858
rect 825 1818 845 1822
rect 914 1801 918 1813
rect 922 1801 926 1813
rect 474 1769 478 1781
rect 483 1769 487 1781
rect 492 1769 496 1781
rect 516 1769 520 1781
rect 524 1769 528 1781
rect 827 1756 831 1796
rect 835 1756 839 1796
rect 714 1727 718 1747
rect 722 1727 726 1747
rect 864 1728 868 1738
rect 872 1728 876 1738
rect 459 1696 463 1708
rect 467 1696 471 1708
rect 498 1680 502 1704
rect 507 1680 511 1704
rect 516 1680 520 1704
rect 526 1674 530 1698
rect 535 1674 539 1698
rect 544 1674 548 1698
rect 459 1641 463 1653
rect 467 1641 471 1653
rect 811 1697 815 1717
rect 819 1697 823 1717
rect 932 1659 936 1671
rect 940 1659 944 1671
rect 971 1643 975 1667
rect 980 1643 984 1667
rect 989 1643 993 1667
rect 999 1637 1003 1661
rect 1008 1637 1012 1661
rect 1017 1637 1021 1661
rect 932 1604 936 1616
rect 940 1604 944 1616
rect 472 1577 476 1589
rect 481 1577 485 1589
rect 490 1577 494 1589
rect 514 1577 518 1589
rect 522 1577 526 1589
rect 827 1588 847 1592
rect 827 1580 847 1584
rect 458 1500 462 1512
rect 466 1500 470 1512
rect 829 1518 833 1558
rect 837 1518 841 1558
rect 497 1484 501 1508
rect 506 1484 510 1508
rect 515 1484 519 1508
rect 525 1478 529 1502
rect 534 1478 538 1502
rect 543 1478 547 1502
rect 733 1490 737 1510
rect 741 1490 745 1510
rect 866 1490 870 1500
rect 874 1490 878 1500
rect 458 1445 462 1457
rect 466 1445 470 1457
rect 813 1459 817 1479
rect 821 1459 825 1479
rect 693 1385 697 1397
rect 701 1385 705 1397
rect 732 1369 736 1393
rect 741 1369 745 1393
rect 750 1369 754 1393
rect 760 1363 764 1387
rect 769 1363 773 1387
rect 778 1363 782 1387
rect 693 1330 697 1342
rect 701 1330 705 1342
<< polysilicon >>
rect 793 2250 796 2252
rect 806 2250 824 2252
rect 844 2250 847 2252
rect 480 2235 482 2238
rect 490 2235 492 2238
rect 522 2235 524 2238
rect 480 2200 482 2223
rect 490 2200 492 2223
rect 522 2205 524 2223
rect 831 2212 833 2215
rect 710 2205 712 2212
rect 717 2205 719 2212
rect 743 2205 745 2212
rect 770 2205 772 2212
rect 793 2205 795 2212
rect 522 2195 524 2198
rect 480 2183 482 2187
rect 490 2183 492 2187
rect 673 2164 675 2167
rect 469 2146 471 2149
rect 508 2142 510 2145
rect 518 2142 520 2145
rect 710 2161 712 2164
rect 717 2161 719 2164
rect 743 2161 745 2165
rect 770 2161 772 2165
rect 793 2161 795 2165
rect 831 2157 833 2172
rect 868 2154 870 2157
rect 469 2120 471 2134
rect 536 2136 538 2139
rect 546 2136 548 2139
rect 469 2111 471 2114
rect 508 2109 510 2118
rect 518 2108 520 2118
rect 673 2126 675 2144
rect 696 2127 698 2134
rect 720 2127 722 2134
rect 741 2127 743 2134
rect 758 2127 760 2134
rect 776 2128 778 2135
rect 815 2133 817 2136
rect 673 2113 675 2116
rect 469 2091 471 2094
rect 469 2065 471 2079
rect 508 2077 510 2104
rect 518 2077 520 2103
rect 536 2101 538 2112
rect 536 2077 538 2097
rect 546 2090 548 2112
rect 868 2129 870 2144
rect 815 2095 817 2113
rect 546 2077 548 2086
rect 696 2083 698 2087
rect 720 2083 722 2087
rect 741 2083 743 2087
rect 758 2083 760 2087
rect 776 2084 778 2088
rect 815 2082 817 2085
rect 508 2062 510 2065
rect 518 2062 520 2065
rect 536 2062 538 2065
rect 546 2062 548 2065
rect 920 2060 922 2063
rect 469 2056 471 2059
rect 959 2056 961 2059
rect 969 2056 971 2059
rect 920 2034 922 2048
rect 987 2050 989 2053
rect 997 2050 999 2053
rect 920 2025 922 2028
rect 959 2023 961 2032
rect 969 2022 971 2032
rect 789 2016 792 2018
rect 802 2016 820 2018
rect 840 2016 843 2018
rect 920 2005 922 2008
rect 471 2000 473 2003
rect 481 2000 483 2003
rect 513 2000 515 2003
rect 827 1990 829 1993
rect 471 1965 473 1988
rect 481 1965 483 1988
rect 513 1970 515 1988
rect 723 1983 725 1990
rect 730 1983 732 1990
rect 756 1983 758 1990
rect 783 1983 785 1990
rect 513 1960 515 1963
rect 471 1948 473 1952
rect 481 1948 483 1952
rect 686 1941 688 1944
rect 920 1979 922 1993
rect 959 1991 961 2018
rect 969 1991 971 2017
rect 987 2015 989 2026
rect 987 1991 989 2011
rect 997 2004 999 2026
rect 997 1991 999 2000
rect 959 1976 961 1979
rect 969 1976 971 1979
rect 987 1976 989 1979
rect 997 1976 999 1979
rect 920 1970 922 1973
rect 723 1939 725 1942
rect 730 1939 732 1942
rect 756 1939 758 1943
rect 783 1939 785 1943
rect 827 1935 829 1950
rect 864 1932 866 1935
rect 467 1911 469 1914
rect 506 1907 508 1910
rect 516 1907 518 1910
rect 467 1885 469 1899
rect 534 1901 536 1904
rect 544 1901 546 1904
rect 686 1903 688 1921
rect 709 1905 711 1912
rect 733 1905 735 1912
rect 754 1905 756 1912
rect 771 1905 773 1912
rect 811 1911 813 1914
rect 467 1876 469 1879
rect 506 1874 508 1883
rect 516 1873 518 1883
rect 686 1890 688 1893
rect 467 1856 469 1859
rect 467 1830 469 1844
rect 506 1842 508 1869
rect 516 1842 518 1868
rect 534 1866 536 1877
rect 534 1842 536 1862
rect 544 1855 546 1877
rect 864 1907 866 1922
rect 811 1873 813 1891
rect 709 1861 711 1865
rect 733 1861 735 1865
rect 754 1861 756 1865
rect 771 1861 773 1865
rect 919 1868 921 1871
rect 811 1860 813 1863
rect 958 1864 960 1867
rect 968 1864 970 1867
rect 544 1842 546 1851
rect 919 1842 921 1856
rect 986 1858 988 1861
rect 996 1858 998 1861
rect 919 1833 921 1836
rect 958 1831 960 1840
rect 506 1827 508 1830
rect 516 1827 518 1830
rect 534 1827 536 1830
rect 544 1827 546 1830
rect 968 1830 970 1840
rect 467 1821 469 1824
rect 794 1823 797 1825
rect 807 1823 825 1825
rect 845 1823 848 1825
rect 919 1813 921 1816
rect 832 1796 834 1799
rect 755 1789 757 1796
rect 762 1789 764 1796
rect 788 1789 790 1796
rect 479 1781 481 1784
rect 489 1781 491 1784
rect 521 1781 523 1784
rect 479 1746 481 1769
rect 489 1746 491 1769
rect 521 1751 523 1769
rect 719 1747 721 1750
rect 919 1787 921 1801
rect 958 1799 960 1826
rect 968 1799 970 1825
rect 986 1823 988 1834
rect 986 1799 988 1819
rect 996 1812 998 1834
rect 996 1799 998 1808
rect 958 1784 960 1787
rect 968 1784 970 1787
rect 986 1784 988 1787
rect 996 1784 998 1787
rect 919 1778 921 1781
rect 521 1741 523 1744
rect 479 1729 481 1733
rect 489 1729 491 1733
rect 755 1745 757 1748
rect 762 1745 764 1748
rect 788 1745 790 1749
rect 832 1741 834 1756
rect 869 1738 871 1741
rect 464 1708 466 1711
rect 719 1709 721 1727
rect 741 1711 743 1718
rect 765 1711 767 1718
rect 786 1711 788 1718
rect 816 1717 818 1720
rect 503 1704 505 1707
rect 513 1704 515 1707
rect 464 1682 466 1696
rect 531 1698 533 1701
rect 541 1698 543 1701
rect 464 1673 466 1676
rect 503 1671 505 1680
rect 513 1670 515 1680
rect 719 1696 721 1699
rect 464 1653 466 1656
rect 464 1627 466 1641
rect 503 1639 505 1666
rect 513 1639 515 1665
rect 531 1663 533 1674
rect 531 1639 533 1659
rect 541 1652 543 1674
rect 869 1713 871 1728
rect 816 1679 818 1697
rect 741 1667 743 1671
rect 765 1667 767 1671
rect 786 1667 788 1671
rect 937 1671 939 1674
rect 816 1666 818 1669
rect 976 1667 978 1670
rect 986 1667 988 1670
rect 541 1639 543 1648
rect 937 1645 939 1659
rect 1004 1661 1006 1664
rect 1014 1661 1016 1664
rect 937 1636 939 1639
rect 976 1634 978 1643
rect 986 1633 988 1643
rect 503 1624 505 1627
rect 513 1624 515 1627
rect 531 1624 533 1627
rect 541 1624 543 1627
rect 464 1618 466 1621
rect 937 1616 939 1619
rect 477 1589 479 1592
rect 487 1589 489 1592
rect 519 1589 521 1592
rect 937 1590 939 1604
rect 976 1602 978 1629
rect 986 1602 988 1628
rect 1004 1626 1006 1637
rect 1004 1602 1006 1622
rect 1014 1615 1016 1637
rect 1014 1602 1016 1611
rect 796 1585 799 1587
rect 809 1585 827 1587
rect 847 1585 850 1587
rect 976 1587 978 1590
rect 986 1587 988 1590
rect 1004 1587 1006 1590
rect 1014 1587 1016 1590
rect 937 1581 939 1584
rect 477 1554 479 1577
rect 487 1554 489 1577
rect 519 1559 521 1577
rect 834 1558 836 1561
rect 519 1549 521 1552
rect 776 1551 778 1558
rect 783 1551 785 1558
rect 477 1537 479 1541
rect 487 1537 489 1541
rect 463 1512 465 1515
rect 502 1508 504 1511
rect 512 1508 514 1511
rect 738 1510 740 1513
rect 463 1486 465 1500
rect 530 1502 532 1505
rect 540 1502 542 1505
rect 463 1477 465 1480
rect 502 1475 504 1484
rect 512 1474 514 1484
rect 776 1507 778 1510
rect 783 1507 785 1510
rect 834 1503 836 1518
rect 871 1500 873 1503
rect 463 1457 465 1460
rect 463 1431 465 1445
rect 502 1443 504 1470
rect 512 1443 514 1469
rect 530 1467 532 1478
rect 530 1443 532 1463
rect 540 1456 542 1478
rect 738 1472 740 1490
rect 762 1473 764 1480
rect 786 1473 788 1480
rect 818 1479 820 1482
rect 738 1459 740 1462
rect 540 1443 542 1452
rect 871 1475 873 1490
rect 818 1441 820 1459
rect 502 1428 504 1431
rect 512 1428 514 1431
rect 530 1428 532 1431
rect 540 1428 542 1431
rect 762 1429 764 1433
rect 786 1429 788 1433
rect 818 1428 820 1431
rect 463 1422 465 1425
rect 698 1397 700 1400
rect 737 1393 739 1396
rect 747 1393 749 1396
rect 698 1371 700 1385
rect 765 1387 767 1390
rect 775 1387 777 1390
rect 698 1362 700 1365
rect 737 1360 739 1369
rect 747 1359 749 1369
rect 698 1342 700 1345
rect 698 1316 700 1330
rect 737 1328 739 1355
rect 747 1328 749 1354
rect 765 1352 767 1363
rect 765 1328 767 1348
rect 775 1341 777 1363
rect 775 1328 777 1337
rect 737 1313 739 1316
rect 747 1313 749 1316
rect 765 1313 767 1316
rect 775 1313 777 1316
rect 698 1307 700 1310
<< polycontact >>
rect 810 2252 814 2256
rect 476 2210 480 2214
rect 486 2203 490 2207
rect 518 2209 522 2213
rect 706 2208 710 2212
rect 719 2208 723 2212
rect 739 2208 743 2212
rect 766 2208 770 2212
rect 789 2208 793 2212
rect 827 2157 831 2161
rect 465 2123 469 2127
rect 669 2130 673 2134
rect 692 2130 696 2134
rect 716 2130 720 2134
rect 737 2130 741 2134
rect 754 2130 758 2134
rect 772 2131 776 2135
rect 465 2068 469 2072
rect 534 2097 538 2101
rect 545 2086 549 2090
rect 864 2129 868 2133
rect 811 2099 815 2103
rect 916 2037 920 2041
rect 806 2018 810 2022
rect 467 1975 471 1979
rect 477 1968 481 1972
rect 509 1974 513 1978
rect 719 1986 723 1990
rect 732 1986 736 1990
rect 752 1986 756 1990
rect 779 1986 783 1990
rect 916 1982 920 1986
rect 985 2011 989 2015
rect 996 2000 1000 2004
rect 823 1935 827 1939
rect 682 1907 686 1911
rect 463 1888 467 1892
rect 705 1908 709 1912
rect 729 1908 733 1912
rect 750 1908 754 1912
rect 767 1908 771 1912
rect 463 1833 467 1837
rect 532 1862 536 1866
rect 860 1907 864 1911
rect 807 1877 811 1881
rect 543 1851 547 1855
rect 915 1845 919 1849
rect 811 1825 815 1829
rect 751 1792 755 1796
rect 764 1792 768 1796
rect 784 1792 788 1796
rect 475 1756 479 1760
rect 485 1749 489 1753
rect 517 1755 521 1759
rect 915 1790 919 1794
rect 984 1819 988 1823
rect 995 1808 999 1812
rect 828 1741 832 1745
rect 715 1713 719 1717
rect 737 1714 741 1718
rect 761 1714 765 1718
rect 782 1714 786 1718
rect 460 1685 464 1689
rect 460 1630 464 1634
rect 529 1659 533 1663
rect 865 1713 869 1717
rect 812 1683 816 1687
rect 540 1648 544 1652
rect 933 1648 937 1652
rect 933 1593 937 1597
rect 813 1587 817 1591
rect 1002 1622 1006 1626
rect 1013 1611 1017 1615
rect 473 1564 477 1568
rect 483 1557 487 1561
rect 515 1563 519 1567
rect 772 1554 776 1558
rect 785 1554 789 1558
rect 459 1489 463 1493
rect 830 1503 834 1507
rect 459 1434 463 1438
rect 528 1463 532 1467
rect 734 1476 738 1480
rect 758 1476 762 1480
rect 782 1476 786 1480
rect 539 1452 543 1456
rect 867 1475 871 1479
rect 814 1445 818 1449
rect 694 1374 698 1378
rect 694 1319 698 1323
rect 763 1348 767 1352
rect 774 1337 778 1341
<< metal1 >>
rect 580 2246 583 2279
rect 467 2241 538 2244
rect 475 2235 479 2241
rect 493 2235 497 2241
rect 517 2235 520 2241
rect 484 2220 487 2223
rect 484 2217 497 2220
rect 437 2210 476 2214
rect 494 2213 497 2217
rect 526 2213 529 2223
rect 437 2209 464 2210
rect 494 2209 518 2213
rect 526 2210 575 2213
rect 471 2206 486 2207
rect 437 2203 486 2206
rect 494 2200 497 2209
rect 526 2205 529 2210
rect 475 2181 478 2187
rect 517 2181 520 2198
rect 467 2178 520 2181
rect 463 2152 491 2155
rect 464 2146 467 2152
rect 488 2151 491 2152
rect 488 2148 559 2151
rect 437 2125 447 2127
rect 437 2122 450 2125
rect 455 2123 465 2126
rect 473 2126 476 2134
rect 503 2142 506 2148
rect 522 2142 525 2148
rect 473 2123 494 2126
rect 473 2120 476 2123
rect 464 2110 467 2114
rect 458 2108 482 2110
rect 458 2107 476 2108
rect 481 2107 482 2108
rect 491 2100 494 2123
rect 532 2142 552 2145
rect 532 2136 535 2142
rect 549 2136 552 2142
rect 513 2115 516 2118
rect 513 2112 531 2115
rect 541 2105 544 2112
rect 541 2102 558 2105
rect 463 2099 482 2100
rect 458 2097 482 2099
rect 491 2097 534 2100
rect 464 2091 467 2097
rect 555 2092 558 2102
rect 520 2086 545 2089
rect 520 2084 523 2086
rect 437 2068 450 2071
rect 455 2068 465 2071
rect 473 2071 476 2079
rect 485 2081 523 2084
rect 555 2083 558 2087
rect 485 2071 488 2081
rect 526 2080 558 2083
rect 526 2077 529 2080
rect 473 2068 488 2071
rect 473 2065 476 2068
rect 525 2074 531 2077
rect 464 2055 467 2059
rect 485 2058 490 2061
rect 503 2061 506 2065
rect 550 2061 553 2065
rect 495 2058 559 2061
rect 485 2055 488 2058
rect 458 2052 488 2055
rect 572 2047 575 2210
rect 580 2093 583 2241
rect 596 2237 600 2280
rect 580 2036 583 2087
rect 588 2056 591 2181
rect 458 2006 529 2009
rect 466 2000 470 2006
rect 484 2000 488 2006
rect 508 2000 511 2006
rect 475 1985 478 1988
rect 475 1982 488 1985
rect 441 1975 467 1979
rect 485 1978 488 1982
rect 517 1978 520 1988
rect 588 1978 591 2051
rect 596 2017 600 2232
rect 612 2227 616 2279
rect 605 2065 608 2182
rect 485 1974 509 1978
rect 517 1975 591 1978
rect 441 1968 477 1972
rect 485 1965 488 1974
rect 517 1970 520 1975
rect 466 1946 469 1952
rect 508 1946 511 1963
rect 458 1943 511 1946
rect 461 1917 489 1920
rect 462 1911 465 1917
rect 486 1916 489 1917
rect 486 1913 557 1916
rect 441 1890 444 1891
rect 441 1887 448 1890
rect 441 1886 444 1887
rect 453 1888 463 1891
rect 471 1891 474 1899
rect 501 1907 504 1913
rect 520 1907 523 1913
rect 471 1888 492 1891
rect 471 1885 474 1888
rect 462 1875 465 1879
rect 456 1873 480 1875
rect 456 1872 474 1873
rect 479 1872 480 1873
rect 489 1865 492 1888
rect 530 1907 550 1910
rect 530 1901 533 1907
rect 547 1901 550 1907
rect 511 1880 514 1883
rect 511 1877 529 1880
rect 539 1870 542 1877
rect 588 1870 591 1975
rect 539 1867 556 1870
rect 461 1864 480 1865
rect 456 1862 480 1864
rect 489 1862 532 1865
rect 462 1856 465 1862
rect 553 1856 556 1867
rect 588 1859 591 1865
rect 596 1860 600 2012
rect 605 1930 608 2060
rect 612 2008 616 2221
rect 632 2218 636 2277
rect 621 2074 624 2181
rect 624 2069 625 2074
rect 595 1856 600 1860
rect 518 1851 543 1854
rect 553 1852 601 1856
rect 518 1849 521 1851
rect 441 1832 448 1837
rect 453 1833 463 1836
rect 471 1836 474 1844
rect 483 1846 521 1849
rect 553 1848 556 1852
rect 483 1836 486 1846
rect 524 1845 556 1848
rect 595 1848 599 1852
rect 524 1842 527 1845
rect 471 1833 486 1836
rect 471 1830 474 1833
rect 523 1839 529 1842
rect 595 1841 599 1843
rect 462 1820 465 1824
rect 483 1823 488 1826
rect 501 1826 504 1830
rect 548 1826 551 1830
rect 493 1823 557 1826
rect 483 1820 486 1823
rect 456 1817 486 1820
rect 466 1787 537 1790
rect 474 1781 478 1787
rect 492 1781 496 1787
rect 516 1781 519 1787
rect 605 1772 608 1925
rect 612 1815 616 2003
rect 621 1920 624 2069
rect 632 1998 636 2213
rect 647 2211 652 2278
rect 785 2257 788 2264
rect 785 2254 796 2257
rect 810 2256 814 2264
rect 850 2257 853 2264
rect 844 2254 853 2257
rect 806 2245 824 2248
rect 725 2212 729 2213
rect 703 2211 706 2212
rect 647 2208 706 2211
rect 723 2208 729 2212
rect 736 2208 739 2221
rect 761 2212 764 2232
rect 783 2212 787 2241
rect 811 2236 814 2245
rect 850 2236 853 2254
rect 761 2208 766 2212
rect 783 2208 789 2212
rect 796 2211 800 2212
rect 604 1769 609 1772
rect 483 1766 486 1769
rect 483 1763 496 1766
rect 423 1760 466 1761
rect 423 1756 475 1760
rect 493 1759 496 1763
rect 525 1759 528 1769
rect 605 1759 608 1769
rect 493 1755 517 1759
rect 525 1756 608 1759
rect 432 1749 485 1753
rect 432 1697 436 1749
rect 493 1746 496 1755
rect 525 1751 528 1756
rect 474 1727 477 1733
rect 516 1727 519 1744
rect 605 1734 608 1756
rect 466 1724 519 1727
rect 458 1714 486 1717
rect 459 1708 462 1714
rect 483 1713 486 1714
rect 483 1710 554 1713
rect 432 1696 435 1697
rect 423 1684 445 1687
rect 423 1682 441 1684
rect 450 1685 460 1688
rect 468 1688 471 1696
rect 498 1704 501 1710
rect 517 1704 520 1710
rect 468 1685 489 1688
rect 468 1682 471 1685
rect 423 1681 427 1682
rect 430 1647 435 1674
rect 459 1672 462 1676
rect 453 1670 477 1672
rect 453 1669 471 1670
rect 476 1669 477 1670
rect 486 1662 489 1685
rect 527 1704 547 1707
rect 527 1698 530 1704
rect 544 1698 547 1704
rect 508 1677 511 1680
rect 508 1674 526 1677
rect 536 1667 539 1674
rect 605 1672 608 1729
rect 612 1669 616 1810
rect 621 1726 624 1915
rect 632 1805 636 1993
rect 536 1664 553 1667
rect 458 1661 477 1662
rect 453 1659 477 1661
rect 486 1659 529 1662
rect 423 1642 435 1647
rect 432 1633 435 1642
rect 459 1653 462 1659
rect 550 1653 553 1664
rect 612 1653 615 1669
rect 515 1648 540 1651
rect 550 1650 615 1653
rect 515 1646 518 1648
rect 432 1630 445 1633
rect 450 1630 460 1633
rect 468 1633 471 1641
rect 480 1643 518 1646
rect 550 1645 553 1650
rect 480 1633 483 1643
rect 521 1642 553 1645
rect 612 1642 615 1650
rect 521 1639 524 1642
rect 468 1630 483 1633
rect 468 1627 471 1630
rect 520 1636 526 1639
rect 459 1617 462 1621
rect 480 1620 485 1623
rect 498 1623 501 1627
rect 545 1623 548 1627
rect 490 1620 554 1623
rect 480 1617 483 1620
rect 453 1614 483 1617
rect 464 1595 535 1598
rect 472 1589 476 1595
rect 490 1589 494 1595
rect 514 1589 517 1595
rect 612 1577 615 1637
rect 481 1574 484 1577
rect 481 1571 494 1574
rect 440 1568 466 1569
rect 414 1564 473 1568
rect 491 1567 494 1571
rect 523 1567 526 1577
rect 621 1567 624 1721
rect 414 1563 440 1564
rect 491 1563 515 1567
rect 523 1564 624 1567
rect 632 1567 636 1800
rect 647 1989 652 2208
rect 796 2207 807 2211
rect 796 2205 800 2207
rect 661 2170 689 2173
rect 668 2164 671 2170
rect 705 2155 709 2164
rect 720 2163 725 2164
rect 738 2163 742 2165
rect 720 2158 742 2163
rect 746 2163 750 2165
rect 765 2163 769 2165
rect 746 2158 769 2163
rect 773 2163 777 2165
rect 788 2163 792 2165
rect 773 2158 792 2163
rect 700 2151 718 2155
rect 677 2134 680 2144
rect 661 2130 669 2134
rect 677 2131 692 2134
rect 677 2126 680 2131
rect 689 2130 692 2131
rect 699 2127 703 2136
rect 668 2108 671 2116
rect 661 2105 671 2108
rect 691 2082 695 2087
rect 706 2082 710 2151
rect 713 2130 716 2140
rect 723 2127 727 2158
rect 751 2154 755 2158
rect 778 2155 782 2158
rect 803 2156 807 2207
rect 810 2161 814 2236
rect 819 2218 847 2221
rect 826 2212 829 2218
rect 810 2157 827 2161
rect 835 2160 838 2172
rect 850 2167 891 2170
rect 850 2160 853 2167
rect 856 2160 884 2163
rect 835 2157 853 2160
rect 744 2150 755 2154
rect 761 2151 782 2155
rect 795 2154 807 2156
rect 839 2154 843 2157
rect 795 2152 843 2154
rect 734 2130 737 2140
rect 744 2127 748 2150
rect 751 2130 754 2138
rect 761 2127 765 2151
rect 769 2145 774 2146
rect 769 2131 772 2140
rect 795 2135 799 2152
rect 803 2150 843 2152
rect 863 2154 866 2160
rect 803 2139 831 2142
rect 779 2131 799 2135
rect 779 2128 783 2131
rect 795 2103 799 2131
rect 810 2133 813 2139
rect 834 2130 864 2133
rect 834 2121 837 2130
rect 856 2129 864 2130
rect 872 2132 875 2144
rect 888 2132 891 2167
rect 872 2129 891 2132
rect 833 2117 902 2121
rect 819 2103 822 2113
rect 834 2103 837 2117
rect 795 2099 811 2103
rect 819 2100 837 2103
rect 819 2095 822 2100
rect 715 2082 719 2087
rect 736 2082 740 2087
rect 753 2082 757 2087
rect 771 2082 775 2088
rect 691 2079 775 2082
rect 810 2077 813 2085
rect 799 2074 813 2077
rect 914 2066 942 2069
rect 915 2060 918 2066
rect 939 2065 942 2066
rect 939 2062 1010 2065
rect 888 2038 901 2039
rect 893 2036 901 2038
rect 906 2037 916 2040
rect 924 2040 927 2048
rect 954 2056 957 2062
rect 973 2056 976 2062
rect 924 2037 945 2040
rect 924 2034 927 2037
rect 781 2023 784 2030
rect 781 2020 792 2023
rect 806 2022 810 2030
rect 846 2023 849 2030
rect 915 2024 918 2028
rect 840 2020 849 2023
rect 909 2022 933 2024
rect 909 2021 927 2022
rect 771 2015 772 2017
rect 771 2012 779 2015
rect 753 2003 754 2008
rect 738 1990 742 1993
rect 716 1989 719 1990
rect 647 1986 719 1989
rect 736 1986 742 1990
rect 749 1986 752 2003
rect 776 1986 779 2012
rect 802 2011 820 2014
rect 807 2002 810 2011
rect 846 2002 849 2020
rect 932 2021 933 2022
rect 942 2014 945 2037
rect 983 2056 1003 2059
rect 983 2050 986 2056
rect 1000 2050 1003 2056
rect 964 2029 967 2032
rect 964 2026 982 2029
rect 992 2019 995 2026
rect 992 2016 1009 2019
rect 914 2013 933 2014
rect 909 2011 933 2013
rect 942 2011 985 2014
rect 915 2005 918 2011
rect 1006 2007 1009 2016
rect 647 1795 652 1986
rect 674 1947 702 1950
rect 681 1941 684 1947
rect 718 1933 722 1942
rect 733 1941 738 1942
rect 751 1941 755 1943
rect 733 1936 755 1941
rect 759 1941 763 1943
rect 778 1941 782 1943
rect 759 1936 782 1941
rect 786 1941 790 1943
rect 786 1936 795 1941
rect 717 1929 724 1933
rect 690 1911 693 1921
rect 702 1911 705 1912
rect 674 1907 682 1911
rect 690 1908 705 1911
rect 690 1903 693 1908
rect 712 1905 716 1914
rect 681 1885 684 1893
rect 674 1882 684 1885
rect 704 1860 708 1865
rect 719 1860 723 1929
rect 726 1908 729 1915
rect 736 1905 740 1936
rect 764 1929 768 1936
rect 791 1932 795 1936
rect 806 1939 810 2002
rect 815 1996 843 1999
rect 822 1990 825 1996
rect 971 2000 996 2003
rect 1006 2003 1023 2007
rect 1006 2001 1012 2003
rect 971 1998 974 2000
rect 806 1935 823 1939
rect 831 1938 834 1950
rect 891 1982 901 1985
rect 846 1945 887 1948
rect 846 1938 849 1945
rect 852 1938 880 1941
rect 831 1935 849 1938
rect 835 1932 839 1935
rect 747 1908 750 1925
rect 757 1925 768 1929
rect 774 1928 839 1932
rect 859 1932 862 1938
rect 757 1905 761 1925
rect 764 1908 767 1916
rect 774 1905 778 1928
rect 791 1881 795 1928
rect 799 1917 827 1920
rect 806 1911 809 1917
rect 815 1881 818 1891
rect 830 1908 860 1911
rect 830 1904 833 1908
rect 852 1907 860 1908
rect 868 1910 871 1922
rect 884 1910 887 1945
rect 868 1907 887 1910
rect 891 1904 894 1982
rect 906 1982 916 1985
rect 924 1985 927 1993
rect 936 1995 974 1998
rect 1006 1997 1009 2001
rect 936 1985 939 1995
rect 977 1994 1009 1997
rect 977 1991 980 1994
rect 924 1982 939 1985
rect 924 1979 927 1982
rect 976 1988 982 1991
rect 915 1969 918 1973
rect 936 1972 941 1975
rect 954 1975 957 1979
rect 1001 1975 1004 1979
rect 946 1972 1010 1975
rect 936 1969 939 1972
rect 909 1966 939 1969
rect 830 1901 894 1904
rect 830 1881 833 1901
rect 791 1877 807 1881
rect 815 1878 833 1881
rect 815 1873 818 1878
rect 913 1874 941 1877
rect 728 1860 732 1865
rect 749 1860 753 1865
rect 766 1860 770 1865
rect 914 1868 917 1874
rect 938 1873 941 1874
rect 938 1870 1009 1873
rect 704 1857 771 1860
rect 806 1855 809 1863
rect 795 1852 809 1855
rect 895 1844 900 1847
rect 905 1845 915 1848
rect 923 1848 926 1856
rect 953 1864 956 1870
rect 972 1864 975 1870
rect 923 1845 944 1848
rect 923 1842 926 1845
rect 786 1830 789 1837
rect 786 1827 797 1830
rect 811 1829 815 1837
rect 851 1830 854 1837
rect 914 1832 917 1836
rect 845 1827 854 1830
rect 908 1830 932 1832
rect 908 1829 926 1830
rect 807 1818 825 1821
rect 781 1810 782 1815
rect 812 1810 815 1818
rect 770 1796 774 1800
rect 748 1795 751 1796
rect 647 1792 751 1795
rect 768 1792 774 1796
rect 781 1792 784 1810
rect 414 1552 419 1563
rect 446 1557 483 1561
rect 446 1555 450 1557
rect 408 1547 419 1552
rect 429 1551 450 1555
rect 491 1554 494 1563
rect 523 1559 526 1564
rect 413 1491 418 1547
rect 429 1503 433 1551
rect 472 1535 475 1541
rect 514 1535 517 1552
rect 464 1532 517 1535
rect 457 1518 485 1521
rect 458 1512 461 1518
rect 482 1517 485 1518
rect 482 1514 553 1517
rect 429 1501 435 1503
rect 423 1491 441 1492
rect 413 1488 444 1491
rect 413 1487 441 1488
rect 449 1489 459 1492
rect 467 1492 470 1500
rect 497 1508 500 1514
rect 516 1508 519 1514
rect 467 1489 488 1492
rect 413 1486 425 1487
rect 467 1486 470 1489
rect 431 1454 436 1479
rect 458 1476 461 1480
rect 452 1474 476 1476
rect 452 1473 470 1474
rect 475 1473 476 1474
rect 485 1466 488 1489
rect 526 1508 546 1511
rect 526 1502 529 1508
rect 543 1502 546 1508
rect 507 1481 510 1484
rect 507 1478 525 1481
rect 620 1488 623 1564
rect 535 1471 538 1478
rect 535 1468 552 1471
rect 457 1465 476 1466
rect 452 1463 476 1465
rect 485 1463 528 1466
rect 408 1449 436 1454
rect 431 1438 436 1449
rect 458 1457 461 1463
rect 549 1457 552 1468
rect 620 1461 623 1483
rect 632 1457 636 1562
rect 514 1452 539 1455
rect 549 1453 636 1457
rect 514 1450 517 1452
rect 431 1437 441 1438
rect 431 1434 444 1437
rect 431 1433 441 1434
rect 449 1434 459 1437
rect 467 1437 470 1445
rect 479 1447 517 1450
rect 549 1449 552 1453
rect 479 1437 482 1447
rect 520 1446 552 1449
rect 520 1443 523 1446
rect 467 1434 482 1437
rect 467 1431 470 1434
rect 519 1440 525 1443
rect 458 1421 461 1425
rect 479 1424 484 1427
rect 497 1427 500 1431
rect 544 1427 547 1431
rect 489 1424 553 1427
rect 479 1421 482 1424
rect 452 1418 482 1421
rect 632 1377 636 1453
rect 647 1558 652 1792
rect 707 1753 735 1756
rect 714 1747 717 1753
rect 750 1735 754 1748
rect 765 1747 770 1748
rect 783 1747 787 1749
rect 765 1742 787 1747
rect 791 1747 795 1749
rect 791 1745 797 1747
rect 811 1745 815 1810
rect 851 1809 854 1827
rect 931 1829 932 1830
rect 941 1822 944 1845
rect 982 1864 1002 1867
rect 982 1858 985 1864
rect 999 1858 1002 1864
rect 963 1837 966 1840
rect 963 1834 981 1837
rect 991 1827 994 1834
rect 991 1824 1008 1827
rect 913 1821 932 1822
rect 908 1819 932 1821
rect 941 1819 984 1822
rect 914 1813 917 1819
rect 1005 1816 1008 1824
rect 820 1802 848 1805
rect 827 1796 830 1802
rect 1005 1812 1023 1816
rect 970 1808 995 1811
rect 970 1806 973 1808
rect 791 1742 799 1745
rect 723 1717 726 1727
rect 735 1717 737 1718
rect 707 1713 715 1717
rect 723 1714 737 1717
rect 723 1709 726 1714
rect 744 1711 748 1720
rect 714 1691 717 1699
rect 707 1688 717 1691
rect 736 1666 740 1671
rect 751 1666 755 1735
rect 758 1714 761 1721
rect 768 1711 772 1742
rect 795 1738 799 1742
rect 811 1741 828 1745
rect 836 1744 839 1756
rect 851 1751 892 1754
rect 851 1744 854 1751
rect 857 1744 885 1747
rect 836 1741 854 1744
rect 840 1738 844 1741
rect 795 1735 844 1738
rect 779 1714 782 1730
rect 789 1734 844 1735
rect 864 1738 867 1744
rect 789 1731 802 1734
rect 789 1711 793 1731
rect 796 1687 800 1731
rect 804 1723 832 1726
rect 811 1717 814 1723
rect 820 1687 823 1697
rect 835 1714 865 1717
rect 835 1699 838 1714
rect 857 1713 865 1714
rect 873 1716 876 1728
rect 889 1716 892 1751
rect 873 1713 892 1716
rect 897 1699 900 1793
rect 905 1790 915 1793
rect 923 1793 926 1801
rect 935 1803 973 1806
rect 1005 1805 1008 1812
rect 935 1793 938 1803
rect 976 1802 1008 1805
rect 976 1799 979 1802
rect 923 1790 938 1793
rect 923 1787 926 1790
rect 975 1796 981 1799
rect 914 1777 917 1781
rect 935 1780 940 1783
rect 953 1783 956 1787
rect 1000 1783 1003 1787
rect 945 1780 1009 1783
rect 935 1777 938 1780
rect 908 1774 938 1777
rect 835 1696 900 1699
rect 835 1687 838 1696
rect 796 1683 812 1687
rect 820 1684 838 1687
rect 820 1679 823 1684
rect 760 1666 764 1671
rect 781 1666 785 1671
rect 931 1677 959 1680
rect 932 1671 935 1677
rect 956 1676 959 1677
rect 956 1673 1027 1676
rect 736 1663 795 1666
rect 811 1661 814 1669
rect 800 1658 814 1661
rect 908 1647 918 1650
rect 923 1648 933 1651
rect 941 1651 944 1659
rect 971 1667 974 1673
rect 990 1667 993 1673
rect 941 1648 962 1651
rect 941 1645 944 1648
rect 932 1635 935 1639
rect 926 1633 950 1635
rect 926 1632 944 1633
rect 949 1632 950 1633
rect 959 1625 962 1648
rect 1000 1667 1020 1670
rect 1000 1661 1003 1667
rect 1017 1661 1020 1667
rect 981 1640 984 1643
rect 981 1637 999 1640
rect 1009 1630 1012 1637
rect 1009 1627 1026 1630
rect 931 1624 950 1625
rect 926 1622 950 1624
rect 959 1622 1002 1625
rect 1023 1622 1026 1627
rect 932 1616 935 1622
rect 1023 1618 1041 1622
rect 988 1611 1013 1614
rect 988 1609 991 1611
rect 788 1592 791 1599
rect 788 1589 799 1592
rect 813 1591 817 1599
rect 853 1592 856 1599
rect 847 1589 856 1592
rect 809 1580 827 1583
rect 814 1571 817 1580
rect 853 1571 856 1589
rect 899 1593 918 1596
rect 791 1558 796 1562
rect 647 1555 772 1558
rect 647 1387 652 1555
rect 769 1554 772 1555
rect 789 1554 796 1558
rect 726 1516 754 1519
rect 733 1510 736 1516
rect 771 1501 775 1510
rect 786 1509 791 1510
rect 786 1504 792 1509
rect 813 1507 817 1571
rect 822 1564 850 1567
rect 829 1558 832 1564
rect 766 1497 784 1501
rect 789 1500 793 1504
rect 813 1503 830 1507
rect 838 1506 841 1518
rect 853 1513 894 1516
rect 853 1506 856 1513
rect 859 1506 887 1509
rect 838 1503 856 1506
rect 842 1500 846 1503
rect 742 1480 745 1490
rect 754 1480 757 1481
rect 726 1476 734 1480
rect 742 1477 758 1480
rect 742 1472 745 1477
rect 754 1476 758 1477
rect 765 1473 769 1482
rect 733 1454 736 1462
rect 726 1451 736 1454
rect 757 1428 761 1433
rect 772 1428 776 1497
rect 789 1496 846 1500
rect 866 1500 869 1506
rect 779 1476 782 1483
rect 789 1473 793 1496
rect 798 1449 802 1496
rect 806 1485 834 1488
rect 813 1479 816 1485
rect 822 1449 825 1459
rect 837 1476 867 1479
rect 837 1467 840 1476
rect 859 1475 867 1476
rect 875 1478 878 1490
rect 891 1478 894 1513
rect 875 1475 894 1478
rect 899 1467 902 1593
rect 923 1593 933 1596
rect 941 1596 944 1604
rect 953 1606 991 1609
rect 1023 1608 1026 1618
rect 953 1596 956 1606
rect 994 1605 1026 1608
rect 994 1602 997 1605
rect 941 1593 956 1596
rect 941 1590 944 1593
rect 993 1599 999 1602
rect 932 1580 935 1584
rect 953 1583 958 1586
rect 971 1586 974 1590
rect 1018 1586 1021 1590
rect 963 1583 1027 1586
rect 953 1580 956 1583
rect 926 1577 956 1580
rect 837 1464 902 1467
rect 837 1449 840 1464
rect 798 1445 814 1449
rect 822 1446 840 1449
rect 822 1441 825 1446
rect 781 1428 785 1433
rect 757 1425 799 1428
rect 813 1423 816 1431
rect 802 1420 816 1423
rect 692 1403 720 1406
rect 693 1397 696 1403
rect 717 1402 720 1403
rect 717 1399 788 1402
rect 642 1377 659 1378
rect 631 1376 673 1377
rect 631 1373 679 1376
rect 684 1374 694 1377
rect 702 1377 705 1385
rect 732 1393 735 1399
rect 751 1393 754 1399
rect 702 1374 723 1377
rect 702 1371 705 1374
rect 647 1345 651 1365
rect 693 1361 696 1365
rect 687 1359 711 1361
rect 687 1358 705 1359
rect 710 1358 711 1359
rect 720 1351 723 1374
rect 761 1393 781 1396
rect 761 1387 764 1393
rect 778 1387 781 1393
rect 742 1366 745 1369
rect 742 1363 760 1366
rect 770 1356 773 1363
rect 770 1353 787 1356
rect 692 1350 711 1351
rect 687 1348 711 1350
rect 720 1348 763 1351
rect 784 1350 794 1353
rect 625 1341 669 1345
rect 665 1322 669 1341
rect 693 1342 696 1348
rect 784 1342 787 1350
rect 749 1337 774 1340
rect 784 1338 790 1342
rect 749 1335 752 1337
rect 665 1319 679 1322
rect 684 1319 694 1322
rect 702 1322 705 1330
rect 714 1332 752 1335
rect 784 1334 787 1338
rect 714 1322 717 1332
rect 755 1331 787 1334
rect 755 1328 758 1331
rect 702 1319 717 1322
rect 702 1316 705 1319
rect 754 1325 760 1328
rect 693 1306 696 1310
rect 714 1309 719 1312
rect 732 1312 735 1316
rect 779 1312 782 1316
rect 724 1309 788 1312
rect 714 1306 717 1309
rect 687 1303 717 1306
<< m2contact >>
rect 579 2241 584 2246
rect 450 2121 455 2126
rect 555 2087 560 2092
rect 450 2067 455 2072
rect 595 2232 600 2237
rect 579 2087 584 2093
rect 571 2042 576 2047
rect 587 2051 592 2056
rect 578 2030 583 2036
rect 612 2221 617 2227
rect 604 2060 609 2065
rect 595 2012 600 2017
rect 448 1886 453 1891
rect 588 1865 593 1870
rect 632 2213 637 2218
rect 619 2069 624 2074
rect 611 2003 616 2008
rect 604 1925 609 1930
rect 448 1832 453 1837
rect 595 1843 600 1848
rect 782 2241 787 2246
rect 760 2232 765 2237
rect 735 2221 740 2227
rect 725 2213 730 2218
rect 632 1993 637 1998
rect 621 1915 626 1920
rect 612 1810 617 1815
rect 603 1729 608 1734
rect 430 1691 435 1696
rect 445 1683 450 1688
rect 430 1674 435 1679
rect 631 1800 636 1805
rect 621 1721 626 1726
rect 445 1629 450 1634
rect 610 1637 615 1642
rect 713 2140 718 2145
rect 732 2140 737 2145
rect 751 2138 756 2143
rect 769 2140 774 2145
rect 888 2033 893 2038
rect 901 2035 906 2040
rect 766 2012 771 2017
rect 748 2003 753 2008
rect 737 1993 742 1998
rect 726 1915 731 1920
rect 745 1925 750 1930
rect 764 1916 769 1921
rect 901 1981 906 1986
rect 890 1842 895 1847
rect 900 1843 905 1848
rect 782 1810 787 1815
rect 769 1800 774 1805
rect 430 1496 435 1501
rect 444 1487 449 1492
rect 430 1479 435 1484
rect 632 1562 637 1567
rect 619 1483 624 1488
rect 444 1433 449 1438
rect 758 1721 763 1726
rect 777 1730 782 1735
rect 900 1789 905 1794
rect 903 1645 908 1650
rect 918 1646 923 1651
rect 791 1562 796 1567
rect 779 1483 784 1488
rect 918 1592 923 1597
rect 647 1382 652 1387
rect 679 1372 684 1377
rect 647 1365 652 1370
rect 679 1318 684 1323
<< pm12contact >>
rect 506 2104 511 2109
rect 515 2103 520 2108
rect 504 1869 509 1874
rect 513 1868 518 1873
rect 501 1666 506 1671
rect 510 1665 515 1670
rect 957 2018 962 2023
rect 966 2017 971 2022
rect 500 1470 505 1475
rect 509 1469 514 1474
rect 956 1826 961 1831
rect 965 1825 970 1830
rect 974 1629 979 1634
rect 983 1628 988 1633
rect 735 1355 740 1360
rect 744 1354 749 1359
<< metal2 >>
rect 584 2241 782 2246
rect 600 2232 760 2237
rect 617 2222 735 2227
rect 637 2213 725 2217
rect 769 2145 774 2146
rect 451 2115 454 2121
rect 451 2112 488 2115
rect 485 2109 488 2112
rect 485 2106 506 2109
rect 515 2093 518 2103
rect 452 2090 518 2093
rect 452 2072 455 2090
rect 560 2087 579 2092
rect 713 2074 718 2140
rect 624 2069 718 2074
rect 732 2065 737 2140
rect 609 2060 737 2065
rect 751 2056 756 2138
rect 592 2051 756 2056
rect 769 2047 774 2140
rect 576 2042 774 2047
rect 773 2036 888 2038
rect 583 2033 888 2036
rect 583 2031 778 2033
rect 902 2029 905 2035
rect 902 2026 939 2029
rect 936 2023 939 2026
rect 600 2012 766 2017
rect 771 2012 772 2017
rect 936 2020 957 2023
rect 616 2003 748 2008
rect 753 2003 754 2008
rect 966 2007 969 2017
rect 903 2004 969 2007
rect 637 1994 737 1998
rect 903 1986 906 2004
rect 609 1925 745 1930
rect 626 1915 726 1920
rect 449 1880 452 1886
rect 449 1877 486 1880
rect 483 1874 486 1877
rect 483 1871 504 1874
rect 764 1870 769 1916
rect 513 1858 516 1868
rect 593 1865 769 1870
rect 450 1855 516 1858
rect 450 1837 453 1855
rect 600 1843 890 1847
rect 901 1837 904 1843
rect 901 1834 938 1837
rect 935 1831 938 1834
rect 935 1828 956 1831
rect 965 1815 968 1825
rect 617 1810 782 1815
rect 902 1812 968 1815
rect 636 1800 769 1805
rect 902 1794 905 1812
rect 602 1734 777 1735
rect 602 1730 603 1734
rect 608 1730 777 1734
rect 626 1721 758 1726
rect 430 1679 435 1691
rect 446 1677 449 1683
rect 446 1674 483 1677
rect 480 1671 483 1674
rect 480 1668 501 1671
rect 510 1655 513 1665
rect 447 1652 513 1655
rect 447 1634 450 1652
rect 903 1642 908 1645
rect 615 1637 908 1642
rect 919 1640 922 1646
rect 919 1637 956 1640
rect 953 1634 956 1637
rect 953 1631 974 1634
rect 983 1618 986 1628
rect 920 1615 986 1618
rect 920 1597 923 1615
rect 637 1562 791 1567
rect 430 1484 435 1496
rect 445 1481 448 1487
rect 624 1483 779 1488
rect 445 1478 482 1481
rect 479 1475 482 1478
rect 479 1472 500 1475
rect 509 1459 512 1469
rect 446 1456 512 1459
rect 446 1438 449 1456
rect 647 1370 652 1382
rect 680 1366 683 1372
rect 680 1363 717 1366
rect 714 1360 717 1363
rect 714 1357 735 1360
rect 744 1344 747 1354
rect 681 1341 747 1344
rect 681 1323 684 1341
<< m123contact >>
rect 458 2152 463 2157
rect 458 2099 463 2104
rect 476 2103 481 2108
rect 490 2058 495 2063
rect 909 2066 914 2071
rect 909 2013 914 2018
rect 927 2017 932 2022
rect 941 1972 946 1977
rect 456 1917 461 1922
rect 456 1864 461 1869
rect 474 1868 479 1873
rect 908 1874 913 1879
rect 488 1823 493 1828
rect 908 1821 913 1826
rect 926 1825 931 1830
rect 940 1780 945 1785
rect 453 1714 458 1719
rect 926 1677 931 1682
rect 453 1661 458 1666
rect 471 1665 476 1670
rect 485 1620 490 1625
rect 926 1624 931 1629
rect 944 1628 949 1633
rect 958 1583 963 1588
rect 452 1518 457 1523
rect 452 1465 457 1470
rect 470 1469 475 1474
rect 484 1424 489 1429
rect 687 1403 692 1408
rect 687 1350 692 1355
rect 705 1354 710 1359
rect 719 1309 724 1314
<< metal3 >>
rect 458 2104 461 2152
rect 481 2103 493 2106
rect 490 2063 493 2103
rect 909 2018 912 2066
rect 932 2017 944 2020
rect 941 1977 944 2017
rect 456 1869 459 1917
rect 479 1868 491 1871
rect 488 1828 491 1868
rect 908 1826 911 1874
rect 931 1825 943 1828
rect 940 1785 943 1825
rect 453 1666 456 1714
rect 476 1665 488 1668
rect 485 1625 488 1665
rect 926 1629 929 1677
rect 949 1628 961 1631
rect 958 1588 961 1628
rect 452 1470 455 1518
rect 475 1469 487 1472
rect 484 1429 487 1469
rect 687 1355 690 1403
rect 710 1354 722 1357
rect 719 1314 722 1354
<< labels >>
rlabel metal1 476 2052 480 2055 1 gnd
rlabel metal1 526 2058 529 2060 1 gnd
rlabel metal1 474 2108 475 2110 1 gnd
rlabel metal1 470 2152 473 2154 5 vdd
rlabel metal1 471 2098 474 2100 1 vdd
rlabel metal1 447 2122 448 2125 1 a3
rlabel metal1 447 2068 448 2071 1 b3
rlabel m2contact 555 2087 559 2091 7 p3
rlabel metal1 533 2211 534 2212 7 g3
rlabel metal1 470 2205 471 2206 3 b3
rlabel metal1 469 2212 470 2213 3 a3
rlabel metal1 493 2243 493 2243 5 vdd!
rlabel metal1 493 2179 493 2179 1 gnd!
rlabel metal1 484 1944 484 1944 1 gnd!
rlabel metal1 484 2008 484 2008 5 vdd!
rlabel metal1 459 1977 460 1978 3 a2
rlabel metal1 461 1970 462 1971 3 b2
rlabel metal1 524 1976 525 1977 7 g2
rlabel metal1 553 1852 557 1856 1 p2
rlabel metal1 445 1833 446 1836 1 b2
rlabel metal1 445 1887 446 1890 1 a2
rlabel metal1 469 1863 472 1865 1 vdd
rlabel metal1 468 1917 471 1919 5 vdd
rlabel metal1 472 1873 473 1875 1 gnd
rlabel metal1 524 1823 527 1825 1 gnd
rlabel metal1 474 1817 478 1820 1 gnd
rlabel metal1 471 1614 475 1617 1 gnd
rlabel metal1 521 1620 524 1622 1 gnd
rlabel metal1 469 1670 470 1672 1 gnd
rlabel metal1 465 1714 468 1716 5 vdd
rlabel metal1 466 1660 469 1662 1 vdd
rlabel metal1 442 1630 443 1633 1 b1
rlabel metal1 442 1684 443 1687 1 a1
rlabel space 550 1649 554 1653 1 p1
rlabel metal1 492 1725 492 1725 1 gnd!
rlabel metal1 492 1789 492 1789 5 vdd!
rlabel metal1 468 1758 469 1759 3 a1
rlabel metal1 469 1751 470 1752 3 b1
rlabel metal1 532 1757 533 1758 7 g1
rlabel metal1 549 1453 553 1457 7 p0
rlabel metal1 465 1464 468 1466 1 vdd
rlabel metal1 464 1518 467 1520 5 vdd
rlabel metal1 468 1474 469 1476 1 gnd
rlabel metal1 520 1424 523 1426 1 gnd
rlabel metal1 470 1418 474 1421 1 gnd
rlabel metal1 490 1597 490 1597 5 vdd!
rlabel metal1 490 1533 490 1533 1 gnd!
rlabel metal1 465 1566 466 1567 3 a0
rlabel metal1 467 1559 468 1560 3 b0
rlabel metal1 530 1565 531 1566 7 g0
rlabel metal1 787 2209 788 2210 1 p3
rlabel metal1 764 2209 765 2210 1 p2
rlabel metal1 737 2209 738 2210 1 p1
rlabel metal1 770 2132 771 2133 1 g3
rlabel metal1 735 2131 736 2132 1 g1
rlabel metal1 714 2131 715 2132 1 g0
rlabel metal1 803 2075 805 2076 1 gnd
rlabel metal1 811 2140 813 2141 1 vdd
rlabel metal1 725 2209 726 2211 1 p0
rlabel metal1 869 2161 876 2162 1 vdd
rlabel metal1 832 2219 839 2220 1 vdd
rlabel metal1 819 2157 825 2161 1 clk
rlabel metal1 834 2100 837 2133 1 c3
rlabel metal1 796 2207 807 2211 1 c3bar
rlabel metal1 689 2130 692 2134 3 clk
rlabel metal1 699 2127 703 2136 1 gnd
rlabel metal1 677 2131 689 2134 1 clk
rlabel metal1 661 2130 669 2134 1 clk_org
rlabel metal1 661 2106 663 2107 1 gnd
rlabel metal1 669 2171 671 2172 1 vdd
rlabel metal1 752 2131 753 2132 1 g2
rlabel metal1 811 2236 814 2248 3 clk
rlabel metal1 810 2256 814 2264 3 clk_org
rlabel metal1 786 2262 787 2264 3 gnd
rlabel metal1 851 2254 852 2256 3 vdd
rlabel metal1 847 2020 848 2022 3 vdd
rlabel metal1 782 2028 783 2030 3 gnd
rlabel metal1 806 2022 810 2030 3 clk_org
rlabel metal1 807 2002 810 2014 3 clk
rlabel metal1 682 1948 684 1949 1 vdd
rlabel metal1 674 1883 676 1884 1 gnd
rlabel metal1 674 1907 682 1911 1 clk_org
rlabel metal1 690 1908 702 1911 1 clk
rlabel metal1 830 1878 833 1911 1 c2
rlabel metal1 791 1877 795 1941 1 c2bar
rlabel metal1 712 1905 716 1914 1 gnd
rlabel metal1 702 1908 705 1912 3 clk
rlabel metal1 738 1987 739 1989 1 p0
rlabel metal1 727 1909 728 1910 1 g0
rlabel metal1 748 1909 749 1910 1 g1
rlabel metal1 765 1909 766 1910 1 g2
rlabel metal1 750 1987 751 1988 1 p1
rlabel metal1 777 1987 778 1988 1 p2
rlabel metal1 815 1935 821 1939 1 clk
rlabel metal1 828 1997 835 1998 1 vdd
rlabel metal1 865 1939 872 1940 1 vdd
rlabel metal1 807 1918 809 1919 1 vdd
rlabel metal1 799 1853 801 1854 1 gnd
rlabel metal1 898 1982 899 1985 1 c2
rlabel metal1 927 1966 931 1969 1 gnd
rlabel metal1 977 1972 980 1974 1 gnd
rlabel metal1 925 2022 926 2024 1 gnd
rlabel metal1 921 2066 924 2068 5 vdd
rlabel metal1 922 2012 925 2014 1 vdd
rlabel metal1 898 2036 899 2039 1 p3
rlabel metal1 715 1754 717 1755 1 vdd
rlabel metal1 707 1689 709 1690 1 gnd
rlabel metal1 707 1713 715 1717 1 clk_org
rlabel metal1 723 1714 735 1717 1 clk
rlabel metal1 812 1809 815 1821 3 clk
rlabel metal1 811 1829 815 1837 3 clk_org
rlabel metal1 787 1835 788 1837 3 gnd
rlabel metal1 852 1827 853 1829 3 vdd
rlabel metal1 835 1684 838 1717 1 c1
rlabel metal1 795 1731 802 1738 1 c1bar
rlabel metal1 782 1793 783 1794 1 p1
rlabel metal1 780 1715 781 1716 1 g1
rlabel metal1 759 1715 760 1716 1 g0
rlabel metal1 770 1793 771 1795 1 p0
rlabel space 734 1714 737 1718 3 clk
rlabel metal1 744 1711 748 1720 1 gnd
rlabel metal1 820 1741 826 1745 1 clk
rlabel metal1 833 1803 840 1804 1 vdd
rlabel metal1 870 1745 877 1746 1 vdd
rlabel metal1 812 1724 814 1725 1 vdd
rlabel metal1 804 1659 806 1660 1 gnd
rlabel metal1 742 1477 754 1480 1 clk
rlabel metal1 726 1476 734 1480 1 clk_org
rlabel metal1 726 1452 728 1453 1 gnd
rlabel metal1 734 1517 736 1518 1 vdd
rlabel metal1 854 1589 855 1591 3 vdd
rlabel metal1 789 1597 790 1599 3 gnd
rlabel metal1 813 1591 817 1599 3 clk_org
rlabel metal1 814 1571 817 1583 3 clk
rlabel metal1 837 1446 840 1479 1 c0
rlabel metal1 789 1496 846 1500 1 c0bar
rlabel metal1 780 1477 781 1478 1 g0
rlabel metal1 791 1555 792 1557 1 p0
rlabel metal1 755 1476 758 1480 3 clk
rlabel metal1 765 1473 769 1482 1 gnd
rlabel metal1 822 1503 828 1507 1 clk
rlabel metal1 835 1565 842 1566 1 vdd
rlabel metal1 872 1507 879 1508 1 vdd
rlabel metal1 814 1486 816 1487 1 vdd
rlabel metal1 806 1421 808 1422 1 gnd
rlabel metal1 901 2119 901 2119 1 c3
rlabel metal1 897 1790 898 1793 1 c1
rlabel metal1 897 1844 898 1847 1 p2
rlabel metal1 921 1820 924 1822 1 vdd
rlabel metal1 920 1874 923 1876 5 vdd
rlabel metal1 924 1830 925 1832 1 gnd
rlabel metal1 976 1780 979 1782 1 gnd
rlabel metal1 926 1774 930 1777 1 gnd
rlabel metal1 788 1340 788 1340 1 s0in
rlabel metal1 676 1373 677 1376 1 p0
rlabel metal1 700 1349 703 1351 1 vdd
rlabel metal1 699 1403 702 1405 5 vdd
rlabel metal1 703 1359 704 1361 1 gnd
rlabel metal1 755 1309 758 1311 1 gnd
rlabel metal1 705 1303 709 1306 1 gnd
rlabel metal1 771 1555 771 1555 1 cin2
rlabel metal1 749 1793 749 1793 1 cin2
rlabel metal1 716 1988 716 1988 1 cin2
rlabel metal1 704 2210 704 2210 1 cin2
rlabel metal1 441 1488 442 1491 1 a0
rlabel metal1 441 1434 442 1437 1 b0
rlabel metal1 915 1593 916 1596 1 c0
rlabel metal1 942 1633 943 1635 1 gnd
rlabel metal1 915 1647 916 1650 1 p1
rlabel metal1 939 1623 942 1625 1 vdd
rlabel metal1 938 1677 941 1679 5 vdd
rlabel metal1 994 1583 997 1585 1 gnd
rlabel metal1 944 1577 948 1580 1 gnd
rlabel metal1 675 1321 675 1321 1 cin
rlabel metal1 1034 1620 1034 1620 1 s1in
rlabel metal1 1017 1814 1017 1814 1 s2in
rlabel metal1 1021 2004 1021 2004 1 s3in
<< end >>
