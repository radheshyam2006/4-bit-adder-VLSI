* SPICE3 file created from D_Flip_Flop.ext - technology: scmos

.option scale=0.09u

M1000 a_n273_n137# a_n280_n116# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=200 ps=120
M1001 a_n273_n137# clk_org a_n269_n105# w_n282_n111# pfet w=25 l=2
+  ad=125 pd=60 as=150 ps=62
M1002 a_n142_n137# a_n187_n105# gnd Gnd nfet w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1003 a_n231_n105# a_n273_n137# a_n237_n137# Gnd nfet w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1004 a_n187_n105# clk_org a_n193_n137# Gnd nfet w=10 l=2
+  ad=50 pd=30 as=60 ps=32
M1005 a_n142_n137# a_n187_n105# vdd w_n155_n111# pfet w=25 l=2
+  ad=125 pd=60 as=500 ps=240
M1006 a_n269_n105# a_n280_n116# vdd w_n282_n111# pfet w=25 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_n193_n137# a_n231_n105# gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_n237_n137# clk_org gnd Gnd nfet w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_n231_n105# clk_org vdd w_n244_n111# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1010 a_n187_n105# a_n231_n105# vdd w_n200_n111# pfet w=25 l=2
+  ad=125 pd=60 as=0 ps=0
C0 a_n187_n105# w_n155_n111# 0.06fF
C1 a_n187_n105# gnd 0.12fF
C2 a_n187_n105# clk_org 0.36fF
C3 a_n269_n105# a_n273_n137# 0.26fF
C4 w_n244_n111# vdd 0.07fF
C5 clk_org a_n280_n116# 0.21fF
C6 a_n269_n105# w_n282_n111# 0.01fF
C7 w_n282_n111# a_n280_n116# 0.06fF
C8 a_n142_n137# a_n187_n105# 0.07fF
C9 w_n200_n111# vdd 0.07fF
C10 w_n244_n111# a_n273_n137# 0.13fF
C11 w_n244_n111# clk_org 0.06fF
C12 w_n244_n111# a_n231_n105# 0.09fF
C13 w_n155_n111# vdd 0.07fF
C14 a_n273_n137# vdd 0.20fF
C15 a_n193_n137# gnd 0.14fF
C16 w_n282_n111# vdd 0.08fF
C17 vdd a_n231_n105# 0.37fF
C18 a_n142_n137# vdd 0.29fF
C19 w_n200_n111# a_n231_n105# 0.06fF
C20 a_n237_n137# gnd 0.14fF
C21 a_n187_n105# vdd 0.37fF
C22 a_n273_n137# gnd 0.24fF
C23 a_n269_n105# vdd 0.29fF
C24 clk_org gnd 0.29fF
C25 a_n142_n137# w_n155_n111# 0.05fF
C26 a_n187_n105# w_n200_n111# 0.09fF
C27 clk_org a_n273_n137# 0.41fF
C28 a_n193_n137# a_n187_n105# 0.10fF
C29 a_n273_n137# w_n282_n111# 0.25fF
C30 gnd a_n231_n105# 0.18fF
C31 a_n237_n137# a_n231_n105# 0.10fF
C32 clk_org w_n282_n111# 0.06fF
C33 a_n142_n137# gnd 0.14fF
C34 a_n273_n137# a_n231_n105# 0.51fF
C35 clk_org a_n231_n105# 0.05fF
C36 a_n193_n137# Gnd 0.01fF
C37 a_n237_n137# Gnd 0.01fF
C38 gnd Gnd 0.08fF
C39 a_n142_n137# Gnd 0.10fF
C40 a_n273_n137# Gnd 0.04fF
C41 vdd Gnd 0.04fF
C42 a_n187_n105# Gnd 0.44fF
C43 a_n231_n105# Gnd 0.48fF
C44 clk_org Gnd 0.44fF
C45 a_n280_n116# Gnd 0.22fF
C46 w_n155_n111# Gnd 0.97fF
C47 w_n200_n111# Gnd 0.97fF
C48 w_n244_n111# Gnd 0.97fF
C49 w_n282_n111# Gnd 0.67fF
