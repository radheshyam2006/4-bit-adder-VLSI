magic
tech scmos
timestamp 1732099764
<< nwell >>
rect 1628 842 1660 879
rect 1666 842 1692 879
rect 1710 842 1736 879
rect 1755 842 1781 879
rect 1853 839 1890 865
rect 1896 839 1924 865
rect 2202 860 2236 888
rect 1844 752 1868 776
rect 1883 766 1917 772
rect 1618 715 1650 752
rect 1656 715 1682 752
rect 1700 715 1726 752
rect 1745 715 1771 752
rect 1883 736 1945 766
rect 2047 760 2075 794
rect 2205 788 2233 842
rect 1911 730 1945 736
rect 2189 729 2217 763
rect 2242 760 2270 784
rect 2289 746 2321 783
rect 2327 746 2353 783
rect 2371 746 2397 783
rect 2416 746 2442 783
rect 2449 743 2477 777
rect 1844 697 1868 721
rect 2295 666 2319 690
rect 2334 680 2368 686
rect 1629 608 1661 645
rect 1667 608 1693 645
rect 1711 608 1737 645
rect 1756 608 1782 645
rect 1844 604 1881 630
rect 1887 604 1915 630
rect 2198 626 2232 654
rect 2334 650 2396 680
rect 2362 644 2396 650
rect 1634 483 1666 520
rect 1672 483 1698 520
rect 1716 483 1742 520
rect 1761 483 1787 520
rect 1842 517 1866 541
rect 2060 537 2088 571
rect 2201 566 2229 620
rect 2295 611 2319 635
rect 2419 632 2451 669
rect 2457 632 2483 669
rect 2501 632 2527 669
rect 2546 632 2572 669
rect 2579 630 2607 664
rect 1881 531 1915 537
rect 1881 501 1943 531
rect 2185 507 2213 541
rect 2238 538 2266 562
rect 1909 495 1943 501
rect 1842 462 1866 486
rect 2294 474 2318 498
rect 2333 488 2367 494
rect 2203 433 2237 461
rect 2333 458 2395 488
rect 2361 452 2395 458
rect 1631 389 1663 426
rect 1669 389 1695 426
rect 1713 389 1739 426
rect 1758 389 1784 426
rect 1852 385 1889 411
rect 1895 385 1923 411
rect 2093 343 2121 377
rect 2206 372 2234 426
rect 2294 419 2318 443
rect 2427 441 2459 478
rect 2465 441 2491 478
rect 2509 441 2535 478
rect 2554 441 2580 478
rect 2586 439 2614 473
rect 1839 314 1863 338
rect 1878 328 1912 334
rect 1642 275 1674 312
rect 1680 275 1706 312
rect 1724 275 1750 312
rect 1769 275 1795 312
rect 1878 298 1940 328
rect 2190 313 2218 347
rect 2243 344 2271 368
rect 1906 292 1940 298
rect 1839 259 1863 283
rect 2312 277 2336 301
rect 2351 291 2385 297
rect 2351 261 2413 291
rect 2379 255 2413 261
rect 2448 247 2480 284
rect 2486 247 2512 284
rect 2530 247 2556 284
rect 2575 247 2601 284
rect 1629 180 1661 217
rect 1667 180 1693 217
rect 1711 180 1737 217
rect 1756 180 1782 217
rect 1850 193 1887 219
rect 1893 193 1921 219
rect 2205 195 2239 223
rect 2312 222 2336 246
rect 2609 245 2637 279
rect 1634 82 1666 119
rect 1672 82 1698 119
rect 1716 82 1742 119
rect 1761 82 1787 119
rect 1838 118 1862 142
rect 1877 132 1911 138
rect 1877 102 1939 132
rect 2112 106 2140 140
rect 2208 134 2236 188
rect 1905 96 1939 102
rect 1838 63 1862 87
rect 2192 75 2220 109
rect 2245 106 2273 130
rect 1773 -25 1805 12
rect 1811 -25 1837 12
rect 1855 -25 1881 12
rect 1900 -25 1926 12
rect 1949 -29 1977 15
rect 1983 -29 2011 20
rect 2073 3 2097 27
rect 2112 17 2146 23
rect 2112 -13 2174 17
rect 2140 -19 2174 -13
rect 2210 -21 2242 16
rect 2248 -21 2274 16
rect 2292 -21 2318 16
rect 2337 -21 2363 16
rect 2371 -23 2399 11
rect 2073 -52 2097 -28
<< ntransistor >>
rect 2182 874 2192 876
rect 1635 816 1637 826
rect 1671 816 1673 826
rect 1679 816 1681 826
rect 1715 816 1717 826
rect 1723 816 1725 826
rect 1766 816 1768 826
rect 1866 811 1868 824
rect 1876 811 1878 824
rect 1908 822 1910 829
rect 2096 788 2098 829
rect 2103 788 2105 829
rect 2129 789 2131 829
rect 2156 789 2158 829
rect 2179 789 2181 829
rect 1855 738 1857 744
rect 2059 740 2061 750
rect 1625 689 1627 699
rect 1661 689 1663 699
rect 1669 689 1671 699
rect 1705 689 1707 699
rect 1713 689 1715 699
rect 1756 689 1758 699
rect 2082 711 2084 751
rect 2106 711 2108 751
rect 2127 711 2129 751
rect 2144 711 2146 751
rect 2162 712 2164 752
rect 2296 720 2298 730
rect 2332 720 2334 730
rect 2340 720 2342 730
rect 2376 720 2378 730
rect 2384 720 2386 730
rect 2427 720 2429 730
rect 2461 723 2463 733
rect 2201 709 2203 719
rect 1894 689 1896 701
rect 1904 689 1906 701
rect 1922 689 1924 701
rect 1932 689 1934 701
rect 1855 683 1857 689
rect 2306 652 2308 658
rect 2178 640 2188 642
rect 1636 582 1638 592
rect 1672 582 1674 592
rect 1680 582 1682 592
rect 1716 582 1718 592
rect 1724 582 1726 592
rect 1767 582 1769 592
rect 1857 576 1859 589
rect 1867 576 1869 589
rect 1899 587 1901 594
rect 2109 566 2111 607
rect 2116 566 2118 607
rect 2142 567 2144 607
rect 2169 567 2171 607
rect 2345 603 2347 615
rect 2355 603 2357 615
rect 2373 603 2375 615
rect 2383 603 2385 615
rect 2426 606 2428 616
rect 2462 606 2464 616
rect 2470 606 2472 616
rect 2506 606 2508 616
rect 2514 606 2516 616
rect 2557 606 2559 616
rect 2591 610 2593 620
rect 2306 597 2308 603
rect 1853 503 1855 509
rect 2072 517 2074 527
rect 1641 457 1643 467
rect 1677 457 1679 467
rect 1685 457 1687 467
rect 1721 457 1723 467
rect 1729 457 1731 467
rect 1772 457 1774 467
rect 2095 489 2097 529
rect 2119 489 2121 529
rect 2140 489 2142 529
rect 2157 489 2159 529
rect 2197 487 2199 497
rect 1892 454 1894 466
rect 1902 454 1904 466
rect 1920 454 1922 466
rect 1930 454 1932 466
rect 2305 460 2307 466
rect 1853 448 1855 454
rect 2183 447 2193 449
rect 1638 363 1640 373
rect 1674 363 1676 373
rect 1682 363 1684 373
rect 1718 363 1720 373
rect 1726 363 1728 373
rect 1769 363 1771 373
rect 1865 357 1867 370
rect 1875 357 1877 370
rect 1907 368 1909 375
rect 2141 372 2143 413
rect 2148 372 2150 413
rect 2174 373 2176 413
rect 2344 411 2346 423
rect 2354 411 2356 423
rect 2372 411 2374 423
rect 2382 411 2384 423
rect 2434 415 2436 425
rect 2470 415 2472 425
rect 2478 415 2480 425
rect 2514 415 2516 425
rect 2522 415 2524 425
rect 2565 415 2567 425
rect 2598 419 2600 429
rect 2305 405 2307 411
rect 1850 300 1852 306
rect 2105 323 2107 333
rect 1649 249 1651 259
rect 1685 249 1687 259
rect 1693 249 1695 259
rect 1729 249 1731 259
rect 1737 249 1739 259
rect 1780 249 1782 259
rect 2127 295 2129 335
rect 2151 295 2153 335
rect 2172 295 2174 335
rect 2202 293 2204 303
rect 2323 263 2325 269
rect 1889 251 1891 263
rect 1899 251 1901 263
rect 1917 251 1919 263
rect 1927 251 1929 263
rect 1850 245 1852 251
rect 2362 214 2364 226
rect 2372 214 2374 226
rect 2390 214 2392 226
rect 2400 214 2402 226
rect 2455 221 2457 231
rect 2491 221 2493 231
rect 2499 221 2501 231
rect 2535 221 2537 231
rect 2543 221 2545 231
rect 2586 221 2588 231
rect 2621 225 2623 235
rect 2185 209 2195 211
rect 2323 208 2325 214
rect 1863 165 1865 178
rect 1873 165 1875 178
rect 1905 176 1907 183
rect 1636 154 1638 164
rect 1672 154 1674 164
rect 1680 154 1682 164
rect 1716 154 1718 164
rect 1724 154 1726 164
rect 1767 154 1769 164
rect 2162 134 2164 175
rect 2169 134 2171 175
rect 1849 104 1851 110
rect 1641 56 1643 66
rect 1677 56 1679 66
rect 1685 56 1687 66
rect 1721 56 1723 66
rect 1729 56 1731 66
rect 1772 56 1774 66
rect 2124 86 2126 96
rect 1888 55 1890 67
rect 1898 55 1900 67
rect 1916 55 1918 67
rect 1926 55 1928 67
rect 2148 57 2150 97
rect 2172 57 2174 97
rect 1849 49 1851 55
rect 2204 55 2206 65
rect 2084 -11 2086 -5
rect 1780 -51 1782 -41
rect 1816 -51 1818 -41
rect 1824 -51 1826 -41
rect 1860 -51 1862 -41
rect 1868 -51 1870 -41
rect 1911 -51 1913 -41
rect 1961 -55 1963 -39
rect 1995 -58 1997 -39
rect 2217 -47 2219 -37
rect 2253 -47 2255 -37
rect 2261 -47 2263 -37
rect 2297 -47 2299 -37
rect 2305 -47 2307 -37
rect 2348 -47 2350 -37
rect 2383 -43 2385 -33
rect 2123 -60 2125 -48
rect 2133 -60 2135 -48
rect 2151 -60 2153 -48
rect 2161 -60 2163 -48
rect 2084 -66 2086 -60
<< ptransistor >>
rect 2210 874 2230 876
rect 1639 848 1641 873
rect 1647 848 1649 873
rect 1677 848 1679 873
rect 1721 848 1723 873
rect 1766 848 1768 873
rect 1866 847 1868 859
rect 1876 847 1878 859
rect 1908 847 1910 859
rect 2217 796 2219 836
rect 1855 758 1857 770
rect 2059 768 2061 788
rect 2254 768 2256 778
rect 1629 721 1631 746
rect 1637 721 1639 746
rect 1667 721 1669 746
rect 1711 721 1713 746
rect 1756 721 1758 746
rect 1894 742 1896 766
rect 1904 742 1906 766
rect 1922 736 1924 760
rect 1932 736 1934 760
rect 1855 703 1857 715
rect 2201 737 2203 757
rect 2300 752 2302 777
rect 2308 752 2310 777
rect 2338 752 2340 777
rect 2382 752 2384 777
rect 2427 752 2429 777
rect 2461 751 2463 771
rect 2306 672 2308 684
rect 2345 656 2347 680
rect 2355 656 2357 680
rect 2373 650 2375 674
rect 2383 650 2385 674
rect 2206 640 2226 642
rect 1640 614 1642 639
rect 1648 614 1650 639
rect 1678 614 1680 639
rect 1722 614 1724 639
rect 1767 614 1769 639
rect 1857 612 1859 624
rect 1867 612 1869 624
rect 1899 612 1901 624
rect 2306 617 2308 629
rect 2213 574 2215 614
rect 2430 638 2432 663
rect 2438 638 2440 663
rect 2468 638 2470 663
rect 2512 638 2514 663
rect 2557 638 2559 663
rect 2591 638 2593 658
rect 2072 545 2074 565
rect 2250 546 2252 556
rect 1853 523 1855 535
rect 1645 489 1647 514
rect 1653 489 1655 514
rect 1683 489 1685 514
rect 1727 489 1729 514
rect 1772 489 1774 514
rect 1892 507 1894 531
rect 1902 507 1904 531
rect 1920 501 1922 525
rect 1930 501 1932 525
rect 1853 468 1855 480
rect 2197 515 2199 535
rect 2305 480 2307 492
rect 2344 464 2346 488
rect 2354 464 2356 488
rect 2372 458 2374 482
rect 2382 458 2384 482
rect 2211 447 2231 449
rect 2305 425 2307 437
rect 1642 395 1644 420
rect 1650 395 1652 420
rect 1680 395 1682 420
rect 1724 395 1726 420
rect 1769 395 1771 420
rect 1865 393 1867 405
rect 1875 393 1877 405
rect 1907 393 1909 405
rect 2218 380 2220 420
rect 2438 447 2440 472
rect 2446 447 2448 472
rect 2476 447 2478 472
rect 2520 447 2522 472
rect 2565 447 2567 472
rect 2598 447 2600 467
rect 2105 351 2107 371
rect 2255 352 2257 362
rect 1850 320 1852 332
rect 1653 281 1655 306
rect 1661 281 1663 306
rect 1691 281 1693 306
rect 1735 281 1737 306
rect 1780 281 1782 306
rect 1889 304 1891 328
rect 1899 304 1901 328
rect 1917 298 1919 322
rect 1927 298 1929 322
rect 1850 265 1852 277
rect 2202 321 2204 341
rect 2323 283 2325 295
rect 2362 267 2364 291
rect 2372 267 2374 291
rect 2390 261 2392 285
rect 2400 261 2402 285
rect 2323 228 2325 240
rect 1640 186 1642 211
rect 1648 186 1650 211
rect 1678 186 1680 211
rect 1722 186 1724 211
rect 1767 186 1769 211
rect 1863 201 1865 213
rect 1873 201 1875 213
rect 1905 201 1907 213
rect 2459 253 2461 278
rect 2467 253 2469 278
rect 2497 253 2499 278
rect 2541 253 2543 278
rect 2586 253 2588 278
rect 2621 253 2623 273
rect 2213 209 2233 211
rect 1849 124 1851 136
rect 2220 142 2222 182
rect 1645 88 1647 113
rect 1653 88 1655 113
rect 1683 88 1685 113
rect 1727 88 1729 113
rect 1772 88 1774 113
rect 1888 108 1890 132
rect 1898 108 1900 132
rect 1916 102 1918 126
rect 1926 102 1928 126
rect 2124 114 2126 134
rect 2257 114 2259 124
rect 1849 69 1851 81
rect 2204 83 2206 103
rect 1784 -19 1786 6
rect 1792 -19 1794 6
rect 1822 -19 1824 6
rect 1866 -19 1868 6
rect 1911 -19 1913 6
rect 1961 -21 1963 9
rect 1995 -21 1997 14
rect 2084 9 2086 21
rect 2123 -7 2125 17
rect 2133 -7 2135 17
rect 2151 -13 2153 11
rect 2161 -13 2163 11
rect 2084 -46 2086 -34
rect 2221 -15 2223 10
rect 2229 -15 2231 10
rect 2259 -15 2261 10
rect 2303 -15 2305 10
rect 2348 -15 2350 10
rect 2383 -15 2385 5
<< ndiffusion >>
rect 2182 876 2192 877
rect 2182 873 2192 874
rect 1634 816 1635 826
rect 1637 816 1638 826
rect 1670 816 1671 826
rect 1673 816 1674 826
rect 1678 816 1679 826
rect 1681 816 1682 826
rect 1714 816 1715 826
rect 1717 816 1718 826
rect 1722 816 1723 826
rect 1725 816 1726 826
rect 1765 816 1766 826
rect 1768 816 1769 826
rect 1865 811 1866 824
rect 1868 811 1876 824
rect 1878 811 1879 824
rect 1907 822 1908 829
rect 1910 822 1911 829
rect 2095 788 2096 829
rect 2098 788 2103 829
rect 2105 788 2106 829
rect 2128 789 2129 829
rect 2131 789 2132 829
rect 2155 789 2156 829
rect 2158 789 2159 829
rect 2178 789 2179 829
rect 2181 789 2182 829
rect 1854 738 1855 744
rect 1857 738 1858 744
rect 2058 740 2059 750
rect 2061 740 2062 750
rect 1624 689 1625 699
rect 1627 689 1628 699
rect 1660 689 1661 699
rect 1663 689 1664 699
rect 1668 689 1669 699
rect 1671 689 1672 699
rect 1704 689 1705 699
rect 1707 689 1708 699
rect 1712 689 1713 699
rect 1715 689 1716 699
rect 1755 689 1756 699
rect 1758 689 1759 699
rect 2081 711 2082 751
rect 2084 711 2085 751
rect 2105 711 2106 751
rect 2108 711 2109 751
rect 2126 711 2127 751
rect 2129 711 2130 751
rect 2143 711 2144 751
rect 2146 711 2147 751
rect 2161 712 2162 752
rect 2164 712 2165 752
rect 2295 720 2296 730
rect 2298 720 2299 730
rect 2331 720 2332 730
rect 2334 720 2335 730
rect 2339 720 2340 730
rect 2342 720 2343 730
rect 2375 720 2376 730
rect 2378 720 2379 730
rect 2383 720 2384 730
rect 2386 720 2387 730
rect 2426 720 2427 730
rect 2429 720 2430 730
rect 2460 723 2461 733
rect 2463 723 2464 733
rect 2200 709 2201 719
rect 2203 709 2204 719
rect 1893 689 1894 701
rect 1896 689 1904 701
rect 1906 689 1907 701
rect 1921 689 1922 701
rect 1924 689 1932 701
rect 1934 689 1935 701
rect 1854 683 1855 689
rect 1857 683 1858 689
rect 2305 652 2306 658
rect 2308 652 2309 658
rect 2178 642 2188 643
rect 2178 639 2188 640
rect 1635 582 1636 592
rect 1638 582 1639 592
rect 1671 582 1672 592
rect 1674 582 1675 592
rect 1679 582 1680 592
rect 1682 582 1683 592
rect 1715 582 1716 592
rect 1718 582 1719 592
rect 1723 582 1724 592
rect 1726 582 1727 592
rect 1766 582 1767 592
rect 1769 582 1770 592
rect 1856 576 1857 589
rect 1859 576 1867 589
rect 1869 576 1870 589
rect 1898 587 1899 594
rect 1901 587 1902 594
rect 2108 566 2109 607
rect 2111 566 2116 607
rect 2118 566 2119 607
rect 2141 567 2142 607
rect 2144 567 2145 607
rect 2168 567 2169 607
rect 2171 567 2172 607
rect 2344 603 2345 615
rect 2347 603 2355 615
rect 2357 603 2358 615
rect 2372 603 2373 615
rect 2375 603 2383 615
rect 2385 603 2386 615
rect 2425 606 2426 616
rect 2428 606 2429 616
rect 2461 606 2462 616
rect 2464 606 2465 616
rect 2469 606 2470 616
rect 2472 606 2473 616
rect 2505 606 2506 616
rect 2508 606 2509 616
rect 2513 606 2514 616
rect 2516 606 2517 616
rect 2556 606 2557 616
rect 2559 606 2560 616
rect 2590 610 2591 620
rect 2593 610 2594 620
rect 2305 597 2306 603
rect 2308 597 2309 603
rect 1852 503 1853 509
rect 1855 503 1856 509
rect 2071 517 2072 527
rect 2074 517 2075 527
rect 1640 457 1641 467
rect 1643 457 1644 467
rect 1676 457 1677 467
rect 1679 457 1680 467
rect 1684 457 1685 467
rect 1687 457 1688 467
rect 1720 457 1721 467
rect 1723 457 1724 467
rect 1728 457 1729 467
rect 1731 457 1732 467
rect 1771 457 1772 467
rect 1774 457 1775 467
rect 2094 489 2095 529
rect 2097 489 2098 529
rect 2118 489 2119 529
rect 2121 489 2122 529
rect 2139 489 2140 529
rect 2142 489 2143 529
rect 2156 489 2157 529
rect 2159 489 2160 529
rect 2196 487 2197 497
rect 2199 487 2200 497
rect 1891 454 1892 466
rect 1894 454 1902 466
rect 1904 454 1905 466
rect 1919 454 1920 466
rect 1922 454 1930 466
rect 1932 454 1933 466
rect 2304 460 2305 466
rect 2307 460 2308 466
rect 1852 448 1853 454
rect 1855 448 1856 454
rect 2183 449 2193 450
rect 2183 446 2193 447
rect 1637 363 1638 373
rect 1640 363 1641 373
rect 1673 363 1674 373
rect 1676 363 1677 373
rect 1681 363 1682 373
rect 1684 363 1685 373
rect 1717 363 1718 373
rect 1720 363 1721 373
rect 1725 363 1726 373
rect 1728 363 1729 373
rect 1768 363 1769 373
rect 1771 363 1772 373
rect 1864 357 1865 370
rect 1867 357 1875 370
rect 1877 357 1878 370
rect 1906 368 1907 375
rect 1909 368 1910 375
rect 2140 372 2141 413
rect 2143 372 2148 413
rect 2150 372 2151 413
rect 2173 373 2174 413
rect 2176 373 2177 413
rect 2343 411 2344 423
rect 2346 411 2354 423
rect 2356 411 2357 423
rect 2371 411 2372 423
rect 2374 411 2382 423
rect 2384 411 2385 423
rect 2433 415 2434 425
rect 2436 415 2437 425
rect 2469 415 2470 425
rect 2472 415 2473 425
rect 2477 415 2478 425
rect 2480 415 2481 425
rect 2513 415 2514 425
rect 2516 415 2517 425
rect 2521 415 2522 425
rect 2524 415 2525 425
rect 2564 415 2565 425
rect 2567 415 2568 425
rect 2597 419 2598 429
rect 2600 419 2601 429
rect 2304 405 2305 411
rect 2307 405 2308 411
rect 1849 300 1850 306
rect 1852 300 1853 306
rect 2104 323 2105 333
rect 2107 323 2108 333
rect 1648 249 1649 259
rect 1651 249 1652 259
rect 1684 249 1685 259
rect 1687 249 1688 259
rect 1692 249 1693 259
rect 1695 249 1696 259
rect 1728 249 1729 259
rect 1731 249 1732 259
rect 1736 249 1737 259
rect 1739 249 1740 259
rect 1779 249 1780 259
rect 1782 249 1783 259
rect 2126 295 2127 335
rect 2129 295 2130 335
rect 2150 295 2151 335
rect 2153 295 2154 335
rect 2171 295 2172 335
rect 2174 295 2175 335
rect 2201 293 2202 303
rect 2204 293 2205 303
rect 2322 263 2323 269
rect 2325 263 2326 269
rect 1888 251 1889 263
rect 1891 251 1899 263
rect 1901 251 1902 263
rect 1916 251 1917 263
rect 1919 251 1927 263
rect 1929 251 1930 263
rect 1849 245 1850 251
rect 1852 245 1853 251
rect 2185 211 2195 212
rect 2361 214 2362 226
rect 2364 214 2372 226
rect 2374 214 2375 226
rect 2389 214 2390 226
rect 2392 214 2400 226
rect 2402 214 2403 226
rect 2454 221 2455 231
rect 2457 221 2458 231
rect 2490 221 2491 231
rect 2493 221 2494 231
rect 2498 221 2499 231
rect 2501 221 2502 231
rect 2534 221 2535 231
rect 2537 221 2538 231
rect 2542 221 2543 231
rect 2545 221 2546 231
rect 2585 221 2586 231
rect 2588 221 2589 231
rect 2620 225 2621 235
rect 2623 225 2624 235
rect 2185 208 2195 209
rect 2322 208 2323 214
rect 2325 208 2326 214
rect 1862 165 1863 178
rect 1865 165 1873 178
rect 1875 165 1876 178
rect 1904 176 1905 183
rect 1907 176 1908 183
rect 1635 154 1636 164
rect 1638 154 1639 164
rect 1671 154 1672 164
rect 1674 154 1675 164
rect 1679 154 1680 164
rect 1682 154 1683 164
rect 1715 154 1716 164
rect 1718 154 1719 164
rect 1723 154 1724 164
rect 1726 154 1727 164
rect 1766 154 1767 164
rect 1769 154 1770 164
rect 2161 134 2162 175
rect 2164 134 2169 175
rect 2171 134 2172 175
rect 1848 104 1849 110
rect 1851 104 1852 110
rect 1640 56 1641 66
rect 1643 56 1644 66
rect 1676 56 1677 66
rect 1679 56 1680 66
rect 1684 56 1685 66
rect 1687 56 1688 66
rect 1720 56 1721 66
rect 1723 56 1724 66
rect 1728 56 1729 66
rect 1731 56 1732 66
rect 1771 56 1772 66
rect 1774 56 1775 66
rect 2123 86 2124 96
rect 2126 86 2127 96
rect 1887 55 1888 67
rect 1890 55 1898 67
rect 1900 55 1901 67
rect 1915 55 1916 67
rect 1918 55 1926 67
rect 1928 55 1929 67
rect 2147 57 2148 97
rect 2150 57 2151 97
rect 2171 57 2172 97
rect 2174 57 2175 97
rect 1848 49 1849 55
rect 1851 49 1852 55
rect 2203 55 2204 65
rect 2206 55 2207 65
rect 2083 -11 2084 -5
rect 2086 -11 2087 -5
rect 1779 -51 1780 -41
rect 1782 -51 1783 -41
rect 1815 -51 1816 -41
rect 1818 -51 1819 -41
rect 1823 -51 1824 -41
rect 1826 -51 1827 -41
rect 1859 -51 1860 -41
rect 1862 -51 1863 -41
rect 1867 -51 1868 -41
rect 1870 -51 1871 -41
rect 1910 -51 1911 -41
rect 1913 -51 1914 -41
rect 1960 -55 1961 -39
rect 1963 -55 1964 -39
rect 1994 -58 1995 -39
rect 1997 -58 1998 -39
rect 2216 -47 2217 -37
rect 2219 -47 2220 -37
rect 2252 -47 2253 -37
rect 2255 -47 2256 -37
rect 2260 -47 2261 -37
rect 2263 -47 2264 -37
rect 2296 -47 2297 -37
rect 2299 -47 2300 -37
rect 2304 -47 2305 -37
rect 2307 -47 2308 -37
rect 2347 -47 2348 -37
rect 2350 -47 2351 -37
rect 2382 -43 2383 -33
rect 2385 -43 2386 -33
rect 2122 -60 2123 -48
rect 2125 -60 2133 -48
rect 2135 -60 2136 -48
rect 2150 -60 2151 -48
rect 2153 -60 2161 -48
rect 2163 -60 2164 -48
rect 2083 -66 2084 -60
rect 2086 -66 2087 -60
<< pdiffusion >>
rect 2210 876 2230 877
rect 1638 848 1639 873
rect 1641 848 1642 873
rect 1646 848 1647 873
rect 1649 848 1650 873
rect 1676 848 1677 873
rect 1679 848 1680 873
rect 1720 848 1721 873
rect 1723 848 1724 873
rect 1765 848 1766 873
rect 1768 848 1769 873
rect 2210 873 2230 874
rect 1865 847 1866 859
rect 1868 847 1870 859
rect 1874 847 1876 859
rect 1878 847 1879 859
rect 1907 847 1908 859
rect 1910 847 1911 859
rect 2216 796 2217 836
rect 2219 796 2220 836
rect 1854 758 1855 770
rect 1857 758 1858 770
rect 2058 768 2059 788
rect 2061 768 2062 788
rect 2253 768 2254 778
rect 2256 768 2257 778
rect 1628 721 1629 746
rect 1631 721 1632 746
rect 1636 721 1637 746
rect 1639 721 1640 746
rect 1666 721 1667 746
rect 1669 721 1670 746
rect 1710 721 1711 746
rect 1713 721 1714 746
rect 1755 721 1756 746
rect 1758 721 1759 746
rect 1893 742 1894 766
rect 1896 742 1898 766
rect 1902 742 1904 766
rect 1906 742 1907 766
rect 1921 736 1922 760
rect 1924 736 1926 760
rect 1930 736 1932 760
rect 1934 736 1935 760
rect 1854 703 1855 715
rect 1857 703 1858 715
rect 2200 737 2201 757
rect 2203 737 2204 757
rect 2299 752 2300 777
rect 2302 752 2303 777
rect 2307 752 2308 777
rect 2310 752 2311 777
rect 2337 752 2338 777
rect 2340 752 2341 777
rect 2381 752 2382 777
rect 2384 752 2385 777
rect 2426 752 2427 777
rect 2429 752 2430 777
rect 2460 751 2461 771
rect 2463 751 2464 771
rect 2305 672 2306 684
rect 2308 672 2309 684
rect 2344 656 2345 680
rect 2347 656 2349 680
rect 2353 656 2355 680
rect 2357 656 2358 680
rect 2206 642 2226 643
rect 2372 650 2373 674
rect 2375 650 2377 674
rect 2381 650 2383 674
rect 2385 650 2386 674
rect 1639 614 1640 639
rect 1642 614 1643 639
rect 1647 614 1648 639
rect 1650 614 1651 639
rect 1677 614 1678 639
rect 1680 614 1681 639
rect 1721 614 1722 639
rect 1724 614 1725 639
rect 1766 614 1767 639
rect 1769 614 1770 639
rect 2206 639 2226 640
rect 1856 612 1857 624
rect 1859 612 1861 624
rect 1865 612 1867 624
rect 1869 612 1870 624
rect 1898 612 1899 624
rect 1901 612 1902 624
rect 2305 617 2306 629
rect 2308 617 2309 629
rect 2212 574 2213 614
rect 2215 574 2216 614
rect 2429 638 2430 663
rect 2432 638 2433 663
rect 2437 638 2438 663
rect 2440 638 2441 663
rect 2467 638 2468 663
rect 2470 638 2471 663
rect 2511 638 2512 663
rect 2514 638 2515 663
rect 2556 638 2557 663
rect 2559 638 2560 663
rect 2590 638 2591 658
rect 2593 638 2594 658
rect 2071 545 2072 565
rect 2074 545 2075 565
rect 2249 546 2250 556
rect 2252 546 2253 556
rect 1852 523 1853 535
rect 1855 523 1856 535
rect 1644 489 1645 514
rect 1647 489 1648 514
rect 1652 489 1653 514
rect 1655 489 1656 514
rect 1682 489 1683 514
rect 1685 489 1686 514
rect 1726 489 1727 514
rect 1729 489 1730 514
rect 1771 489 1772 514
rect 1774 489 1775 514
rect 1891 507 1892 531
rect 1894 507 1896 531
rect 1900 507 1902 531
rect 1904 507 1905 531
rect 1919 501 1920 525
rect 1922 501 1924 525
rect 1928 501 1930 525
rect 1932 501 1933 525
rect 1852 468 1853 480
rect 1855 468 1856 480
rect 2196 515 2197 535
rect 2199 515 2200 535
rect 2304 480 2305 492
rect 2307 480 2308 492
rect 2343 464 2344 488
rect 2346 464 2348 488
rect 2352 464 2354 488
rect 2356 464 2357 488
rect 2371 458 2372 482
rect 2374 458 2376 482
rect 2380 458 2382 482
rect 2384 458 2385 482
rect 2211 449 2231 450
rect 2211 446 2231 447
rect 2304 425 2305 437
rect 2307 425 2308 437
rect 1641 395 1642 420
rect 1644 395 1645 420
rect 1649 395 1650 420
rect 1652 395 1653 420
rect 1679 395 1680 420
rect 1682 395 1683 420
rect 1723 395 1724 420
rect 1726 395 1727 420
rect 1768 395 1769 420
rect 1771 395 1772 420
rect 1864 393 1865 405
rect 1867 393 1869 405
rect 1873 393 1875 405
rect 1877 393 1878 405
rect 1906 393 1907 405
rect 1909 393 1910 405
rect 2217 380 2218 420
rect 2220 380 2221 420
rect 2437 447 2438 472
rect 2440 447 2441 472
rect 2445 447 2446 472
rect 2448 447 2449 472
rect 2475 447 2476 472
rect 2478 447 2479 472
rect 2519 447 2520 472
rect 2522 447 2523 472
rect 2564 447 2565 472
rect 2567 447 2568 472
rect 2597 447 2598 467
rect 2600 447 2601 467
rect 2104 351 2105 371
rect 2107 351 2108 371
rect 2254 352 2255 362
rect 2257 352 2258 362
rect 1849 320 1850 332
rect 1852 320 1853 332
rect 1652 281 1653 306
rect 1655 281 1656 306
rect 1660 281 1661 306
rect 1663 281 1664 306
rect 1690 281 1691 306
rect 1693 281 1694 306
rect 1734 281 1735 306
rect 1737 281 1738 306
rect 1779 281 1780 306
rect 1782 281 1783 306
rect 1888 304 1889 328
rect 1891 304 1893 328
rect 1897 304 1899 328
rect 1901 304 1902 328
rect 1916 298 1917 322
rect 1919 298 1921 322
rect 1925 298 1927 322
rect 1929 298 1930 322
rect 1849 265 1850 277
rect 1852 265 1853 277
rect 2201 321 2202 341
rect 2204 321 2205 341
rect 2322 283 2323 295
rect 2325 283 2326 295
rect 2361 267 2362 291
rect 2364 267 2366 291
rect 2370 267 2372 291
rect 2374 267 2375 291
rect 2389 261 2390 285
rect 2392 261 2394 285
rect 2398 261 2400 285
rect 2402 261 2403 285
rect 2322 228 2323 240
rect 2325 228 2326 240
rect 1639 186 1640 211
rect 1642 186 1643 211
rect 1647 186 1648 211
rect 1650 186 1651 211
rect 1677 186 1678 211
rect 1680 186 1681 211
rect 1721 186 1722 211
rect 1724 186 1725 211
rect 1766 186 1767 211
rect 1769 186 1770 211
rect 1862 201 1863 213
rect 1865 201 1867 213
rect 1871 201 1873 213
rect 1875 201 1876 213
rect 1904 201 1905 213
rect 1907 201 1908 213
rect 2458 253 2459 278
rect 2461 253 2462 278
rect 2466 253 2467 278
rect 2469 253 2470 278
rect 2496 253 2497 278
rect 2499 253 2500 278
rect 2540 253 2541 278
rect 2543 253 2544 278
rect 2585 253 2586 278
rect 2588 253 2589 278
rect 2620 253 2621 273
rect 2623 253 2624 273
rect 2213 211 2233 212
rect 2213 208 2233 209
rect 1848 124 1849 136
rect 1851 124 1852 136
rect 2219 142 2220 182
rect 2222 142 2223 182
rect 1644 88 1645 113
rect 1647 88 1648 113
rect 1652 88 1653 113
rect 1655 88 1656 113
rect 1682 88 1683 113
rect 1685 88 1686 113
rect 1726 88 1727 113
rect 1729 88 1730 113
rect 1771 88 1772 113
rect 1774 88 1775 113
rect 1887 108 1888 132
rect 1890 108 1892 132
rect 1896 108 1898 132
rect 1900 108 1901 132
rect 1915 102 1916 126
rect 1918 102 1920 126
rect 1924 102 1926 126
rect 1928 102 1929 126
rect 2123 114 2124 134
rect 2126 114 2127 134
rect 2256 114 2257 124
rect 2259 114 2260 124
rect 1848 69 1849 81
rect 1851 69 1852 81
rect 2203 83 2204 103
rect 2206 83 2207 103
rect 1783 -19 1784 6
rect 1786 -19 1787 6
rect 1791 -19 1792 6
rect 1794 -19 1795 6
rect 1821 -19 1822 6
rect 1824 -19 1825 6
rect 1865 -19 1866 6
rect 1868 -19 1869 6
rect 1910 -19 1911 6
rect 1913 -19 1914 6
rect 1960 -21 1961 9
rect 1963 -21 1964 9
rect 1994 -21 1995 14
rect 1997 -21 1998 14
rect 2083 9 2084 21
rect 2086 9 2087 21
rect 2122 -7 2123 17
rect 2125 -7 2127 17
rect 2131 -7 2133 17
rect 2135 -7 2136 17
rect 2150 -13 2151 11
rect 2153 -13 2155 11
rect 2159 -13 2161 11
rect 2163 -13 2164 11
rect 2083 -46 2084 -34
rect 2086 -46 2087 -34
rect 2220 -15 2221 10
rect 2223 -15 2224 10
rect 2228 -15 2229 10
rect 2231 -15 2232 10
rect 2258 -15 2259 10
rect 2261 -15 2262 10
rect 2302 -15 2303 10
rect 2305 -15 2306 10
rect 2347 -15 2348 10
rect 2350 -15 2351 10
rect 2382 -15 2383 5
rect 2385 -15 2386 5
<< ndcontact >>
rect 2182 877 2192 881
rect 2182 869 2192 873
rect 1630 816 1634 826
rect 1638 816 1642 826
rect 1666 816 1670 826
rect 1674 816 1678 826
rect 1682 816 1686 826
rect 1710 816 1714 826
rect 1718 816 1722 826
rect 1726 816 1730 826
rect 1761 816 1765 826
rect 1769 816 1773 826
rect 1861 811 1865 824
rect 1879 811 1883 824
rect 1903 822 1907 829
rect 1911 822 1915 829
rect 2091 788 2095 829
rect 2106 788 2111 829
rect 2124 789 2128 829
rect 2132 789 2136 829
rect 2151 789 2155 829
rect 2159 789 2163 829
rect 2174 789 2178 829
rect 2182 789 2186 829
rect 1850 738 1854 744
rect 1858 738 1862 744
rect 2054 740 2058 750
rect 2062 740 2066 750
rect 1620 689 1624 699
rect 1628 689 1632 699
rect 1656 689 1660 699
rect 1664 689 1668 699
rect 1672 689 1676 699
rect 1700 689 1704 699
rect 1708 689 1712 699
rect 1716 689 1720 699
rect 1751 689 1755 699
rect 1759 689 1763 699
rect 2077 711 2081 751
rect 2085 711 2089 751
rect 2101 711 2105 751
rect 2109 711 2113 751
rect 2122 711 2126 751
rect 2130 711 2134 751
rect 2139 711 2143 751
rect 2147 711 2151 751
rect 2157 712 2161 752
rect 2165 712 2169 752
rect 2291 720 2295 730
rect 2299 720 2303 730
rect 2327 720 2331 730
rect 2335 720 2339 730
rect 2343 720 2347 730
rect 2371 720 2375 730
rect 2379 720 2383 730
rect 2387 720 2391 730
rect 2422 720 2426 730
rect 2430 720 2434 730
rect 2456 723 2460 733
rect 2464 723 2468 733
rect 2196 709 2200 719
rect 2204 709 2208 719
rect 1889 689 1893 701
rect 1907 689 1911 701
rect 1917 689 1921 701
rect 1935 689 1939 701
rect 1850 683 1854 689
rect 1858 683 1862 689
rect 2301 652 2305 658
rect 2309 652 2313 658
rect 2178 643 2188 647
rect 2178 635 2188 639
rect 1631 582 1635 592
rect 1639 582 1643 592
rect 1667 582 1671 592
rect 1675 582 1679 592
rect 1683 582 1687 592
rect 1711 582 1715 592
rect 1719 582 1723 592
rect 1727 582 1731 592
rect 1762 582 1766 592
rect 1770 582 1774 592
rect 1852 576 1856 589
rect 1870 576 1874 589
rect 1894 587 1898 594
rect 1902 587 1906 594
rect 2104 566 2108 607
rect 2119 566 2124 607
rect 2137 567 2141 607
rect 2145 567 2149 607
rect 2164 567 2168 607
rect 2172 567 2176 607
rect 2340 603 2344 615
rect 2358 603 2362 615
rect 2368 603 2372 615
rect 2386 603 2390 615
rect 2421 606 2425 616
rect 2429 606 2433 616
rect 2457 606 2461 616
rect 2465 606 2469 616
rect 2473 606 2477 616
rect 2501 606 2505 616
rect 2509 606 2513 616
rect 2517 606 2521 616
rect 2552 606 2556 616
rect 2560 606 2564 616
rect 2586 610 2590 620
rect 2594 610 2598 620
rect 2301 597 2305 603
rect 2309 597 2313 603
rect 1848 503 1852 509
rect 1856 503 1860 509
rect 2067 517 2071 527
rect 2075 517 2079 527
rect 1636 457 1640 467
rect 1644 457 1648 467
rect 1672 457 1676 467
rect 1680 457 1684 467
rect 1688 457 1692 467
rect 1716 457 1720 467
rect 1724 457 1728 467
rect 1732 457 1736 467
rect 1767 457 1771 467
rect 1775 457 1779 467
rect 2090 489 2094 529
rect 2098 489 2102 529
rect 2114 489 2118 529
rect 2122 489 2126 529
rect 2135 489 2139 529
rect 2143 489 2147 529
rect 2152 489 2156 529
rect 2160 489 2164 529
rect 2192 487 2196 497
rect 2200 487 2204 497
rect 1887 454 1891 466
rect 1905 454 1909 466
rect 1915 454 1919 466
rect 1933 454 1937 466
rect 2300 460 2304 466
rect 2308 460 2312 466
rect 1848 448 1852 454
rect 1856 448 1860 454
rect 2183 450 2193 454
rect 2183 442 2193 446
rect 1633 363 1637 373
rect 1641 363 1645 373
rect 1669 363 1673 373
rect 1677 363 1681 373
rect 1685 363 1689 373
rect 1713 363 1717 373
rect 1721 363 1725 373
rect 1729 363 1733 373
rect 1764 363 1768 373
rect 1772 363 1776 373
rect 1860 357 1864 370
rect 1878 357 1882 370
rect 1902 368 1906 375
rect 1910 368 1914 375
rect 2136 372 2140 413
rect 2151 372 2156 413
rect 2169 373 2173 413
rect 2177 373 2181 413
rect 2339 411 2343 423
rect 2357 411 2361 423
rect 2367 411 2371 423
rect 2385 411 2389 423
rect 2429 415 2433 425
rect 2437 415 2441 425
rect 2465 415 2469 425
rect 2473 415 2477 425
rect 2481 415 2485 425
rect 2509 415 2513 425
rect 2517 415 2521 425
rect 2525 415 2529 425
rect 2560 415 2564 425
rect 2568 415 2572 425
rect 2593 419 2597 429
rect 2601 419 2605 429
rect 2300 405 2304 411
rect 2308 405 2312 411
rect 1845 300 1849 306
rect 1853 300 1857 306
rect 2100 323 2104 333
rect 2108 323 2112 333
rect 1644 249 1648 259
rect 1652 249 1656 259
rect 1680 249 1684 259
rect 1688 249 1692 259
rect 1696 249 1700 259
rect 1724 249 1728 259
rect 1732 249 1736 259
rect 1740 249 1744 259
rect 1775 249 1779 259
rect 1783 249 1787 259
rect 2122 295 2126 335
rect 2130 295 2134 335
rect 2146 295 2150 335
rect 2154 295 2158 335
rect 2167 295 2171 335
rect 2175 295 2179 335
rect 2197 293 2201 303
rect 2205 293 2209 303
rect 2318 263 2322 269
rect 2326 263 2330 269
rect 1884 251 1888 263
rect 1902 251 1906 263
rect 1912 251 1916 263
rect 1930 251 1934 263
rect 1845 245 1849 251
rect 1853 245 1857 251
rect 2185 212 2195 216
rect 2357 214 2361 226
rect 2375 214 2379 226
rect 2385 214 2389 226
rect 2403 214 2407 226
rect 2450 221 2454 231
rect 2458 221 2462 231
rect 2486 221 2490 231
rect 2494 221 2498 231
rect 2502 221 2506 231
rect 2530 221 2534 231
rect 2538 221 2542 231
rect 2546 221 2550 231
rect 2581 221 2585 231
rect 2589 221 2593 231
rect 2616 225 2620 235
rect 2624 225 2628 235
rect 2185 204 2195 208
rect 2318 208 2322 214
rect 2326 208 2330 214
rect 1858 165 1862 178
rect 1876 165 1880 178
rect 1900 176 1904 183
rect 1908 176 1912 183
rect 1631 154 1635 164
rect 1639 154 1643 164
rect 1667 154 1671 164
rect 1675 154 1679 164
rect 1683 154 1687 164
rect 1711 154 1715 164
rect 1719 154 1723 164
rect 1727 154 1731 164
rect 1762 154 1766 164
rect 1770 154 1774 164
rect 2157 134 2161 175
rect 2172 134 2177 175
rect 1844 104 1848 110
rect 1852 104 1856 110
rect 1636 56 1640 66
rect 1644 56 1648 66
rect 1672 56 1676 66
rect 1680 56 1684 66
rect 1688 56 1692 66
rect 1716 56 1720 66
rect 1724 56 1728 66
rect 1732 56 1736 66
rect 1767 56 1771 66
rect 1775 56 1779 66
rect 2119 86 2123 96
rect 2127 86 2131 96
rect 1883 55 1887 67
rect 1901 55 1905 67
rect 1911 55 1915 67
rect 1929 55 1933 67
rect 2143 57 2147 97
rect 2151 57 2155 97
rect 2167 57 2171 97
rect 2175 57 2179 97
rect 1844 49 1848 55
rect 1852 49 1856 55
rect 2199 55 2203 65
rect 2207 55 2211 65
rect 2079 -11 2083 -5
rect 2087 -11 2091 -5
rect 1775 -51 1779 -41
rect 1783 -51 1787 -41
rect 1811 -51 1815 -41
rect 1819 -51 1823 -41
rect 1827 -51 1831 -41
rect 1855 -51 1859 -41
rect 1863 -51 1867 -41
rect 1871 -51 1875 -41
rect 1906 -51 1910 -41
rect 1914 -51 1918 -41
rect 1956 -55 1960 -39
rect 1964 -55 1968 -39
rect 1990 -58 1994 -39
rect 1998 -58 2002 -39
rect 2212 -47 2216 -37
rect 2220 -47 2224 -37
rect 2248 -47 2252 -37
rect 2256 -47 2260 -37
rect 2264 -47 2268 -37
rect 2292 -47 2296 -37
rect 2300 -47 2304 -37
rect 2308 -47 2312 -37
rect 2343 -47 2347 -37
rect 2351 -47 2355 -37
rect 2378 -43 2382 -33
rect 2386 -43 2390 -33
rect 2118 -60 2122 -48
rect 2136 -60 2140 -48
rect 2146 -60 2150 -48
rect 2164 -60 2168 -48
rect 2079 -66 2083 -60
rect 2087 -66 2091 -60
<< pdcontact >>
rect 2210 877 2230 881
rect 1634 848 1638 873
rect 1642 848 1646 873
rect 1650 848 1654 873
rect 1672 848 1676 873
rect 1680 848 1684 873
rect 1716 848 1720 873
rect 1724 848 1728 873
rect 1761 848 1765 873
rect 1769 848 1773 873
rect 2210 869 2230 873
rect 1861 847 1865 859
rect 1870 847 1874 859
rect 1879 847 1883 859
rect 1903 847 1907 859
rect 1911 847 1915 859
rect 2212 796 2216 836
rect 2220 796 2224 836
rect 1850 758 1854 770
rect 1858 758 1862 770
rect 2054 768 2058 788
rect 2062 768 2066 788
rect 2249 768 2253 778
rect 2257 768 2261 778
rect 1624 721 1628 746
rect 1632 721 1636 746
rect 1640 721 1644 746
rect 1662 721 1666 746
rect 1670 721 1674 746
rect 1706 721 1710 746
rect 1714 721 1718 746
rect 1751 721 1755 746
rect 1759 721 1763 746
rect 1889 742 1893 766
rect 1898 742 1902 766
rect 1907 742 1911 766
rect 1917 736 1921 760
rect 1926 736 1930 760
rect 1935 736 1939 760
rect 1850 703 1854 715
rect 1858 703 1862 715
rect 2196 737 2200 757
rect 2204 737 2208 757
rect 2295 752 2299 777
rect 2303 752 2307 777
rect 2311 752 2315 777
rect 2333 752 2337 777
rect 2341 752 2345 777
rect 2377 752 2381 777
rect 2385 752 2389 777
rect 2422 752 2426 777
rect 2430 752 2434 777
rect 2456 751 2460 771
rect 2464 751 2468 771
rect 2301 672 2305 684
rect 2309 672 2313 684
rect 2340 656 2344 680
rect 2349 656 2353 680
rect 2358 656 2362 680
rect 2206 643 2226 647
rect 2368 650 2372 674
rect 2377 650 2381 674
rect 2386 650 2390 674
rect 1635 614 1639 639
rect 1643 614 1647 639
rect 1651 614 1655 639
rect 1673 614 1677 639
rect 1681 614 1685 639
rect 1717 614 1721 639
rect 1725 614 1729 639
rect 1762 614 1766 639
rect 1770 614 1774 639
rect 2206 635 2226 639
rect 1852 612 1856 624
rect 1861 612 1865 624
rect 1870 612 1874 624
rect 1894 612 1898 624
rect 1902 612 1906 624
rect 2301 617 2305 629
rect 2309 617 2313 629
rect 2208 574 2212 614
rect 2216 574 2220 614
rect 2425 638 2429 663
rect 2433 638 2437 663
rect 2441 638 2445 663
rect 2463 638 2467 663
rect 2471 638 2475 663
rect 2507 638 2511 663
rect 2515 638 2519 663
rect 2552 638 2556 663
rect 2560 638 2564 663
rect 2586 638 2590 658
rect 2594 638 2598 658
rect 2067 545 2071 565
rect 2075 545 2079 565
rect 2245 546 2249 556
rect 2253 546 2257 556
rect 1848 523 1852 535
rect 1856 523 1860 535
rect 1640 489 1644 514
rect 1648 489 1652 514
rect 1656 489 1660 514
rect 1678 489 1682 514
rect 1686 489 1690 514
rect 1722 489 1726 514
rect 1730 489 1734 514
rect 1767 489 1771 514
rect 1775 489 1779 514
rect 1887 507 1891 531
rect 1896 507 1900 531
rect 1905 507 1909 531
rect 1915 501 1919 525
rect 1924 501 1928 525
rect 1933 501 1937 525
rect 1848 468 1852 480
rect 1856 468 1860 480
rect 2192 515 2196 535
rect 2200 515 2204 535
rect 2300 480 2304 492
rect 2308 480 2312 492
rect 2339 464 2343 488
rect 2348 464 2352 488
rect 2357 464 2361 488
rect 2211 450 2231 454
rect 2367 458 2371 482
rect 2376 458 2380 482
rect 2385 458 2389 482
rect 2211 442 2231 446
rect 2300 425 2304 437
rect 2308 425 2312 437
rect 1637 395 1641 420
rect 1645 395 1649 420
rect 1653 395 1657 420
rect 1675 395 1679 420
rect 1683 395 1687 420
rect 1719 395 1723 420
rect 1727 395 1731 420
rect 1764 395 1768 420
rect 1772 395 1776 420
rect 1860 393 1864 405
rect 1869 393 1873 405
rect 1878 393 1882 405
rect 1902 393 1906 405
rect 1910 393 1914 405
rect 2213 380 2217 420
rect 2221 380 2225 420
rect 2433 447 2437 472
rect 2441 447 2445 472
rect 2449 447 2453 472
rect 2471 447 2475 472
rect 2479 447 2483 472
rect 2515 447 2519 472
rect 2523 447 2527 472
rect 2560 447 2564 472
rect 2568 447 2572 472
rect 2593 447 2597 467
rect 2601 447 2605 467
rect 2100 351 2104 371
rect 2108 351 2112 371
rect 2250 352 2254 362
rect 2258 352 2262 362
rect 1845 320 1849 332
rect 1853 320 1857 332
rect 1648 281 1652 306
rect 1656 281 1660 306
rect 1664 281 1668 306
rect 1686 281 1690 306
rect 1694 281 1698 306
rect 1730 281 1734 306
rect 1738 281 1742 306
rect 1775 281 1779 306
rect 1783 281 1787 306
rect 1884 304 1888 328
rect 1893 304 1897 328
rect 1902 304 1906 328
rect 1912 298 1916 322
rect 1921 298 1925 322
rect 1930 298 1934 322
rect 1845 265 1849 277
rect 1853 265 1857 277
rect 2197 321 2201 341
rect 2205 321 2209 341
rect 2318 283 2322 295
rect 2326 283 2330 295
rect 2357 267 2361 291
rect 2366 267 2370 291
rect 2375 267 2379 291
rect 2385 261 2389 285
rect 2394 261 2398 285
rect 2403 261 2407 285
rect 2318 228 2322 240
rect 2326 228 2330 240
rect 1635 186 1639 211
rect 1643 186 1647 211
rect 1651 186 1655 211
rect 1673 186 1677 211
rect 1681 186 1685 211
rect 1717 186 1721 211
rect 1725 186 1729 211
rect 1762 186 1766 211
rect 1770 186 1774 211
rect 1858 201 1862 213
rect 1867 201 1871 213
rect 1876 201 1880 213
rect 1900 201 1904 213
rect 1908 201 1912 213
rect 2213 212 2233 216
rect 2454 253 2458 278
rect 2462 253 2466 278
rect 2470 253 2474 278
rect 2492 253 2496 278
rect 2500 253 2504 278
rect 2536 253 2540 278
rect 2544 253 2548 278
rect 2581 253 2585 278
rect 2589 253 2593 278
rect 2616 253 2620 273
rect 2624 253 2628 273
rect 2213 204 2233 208
rect 1844 124 1848 136
rect 1852 124 1856 136
rect 2215 142 2219 182
rect 2223 142 2227 182
rect 1640 88 1644 113
rect 1648 88 1652 113
rect 1656 88 1660 113
rect 1678 88 1682 113
rect 1686 88 1690 113
rect 1722 88 1726 113
rect 1730 88 1734 113
rect 1767 88 1771 113
rect 1775 88 1779 113
rect 1883 108 1887 132
rect 1892 108 1896 132
rect 1901 108 1905 132
rect 1911 102 1915 126
rect 1920 102 1924 126
rect 1929 102 1933 126
rect 2119 114 2123 134
rect 2127 114 2131 134
rect 2252 114 2256 124
rect 2260 114 2264 124
rect 1844 69 1848 81
rect 1852 69 1856 81
rect 2199 83 2203 103
rect 2207 83 2211 103
rect 1779 -19 1783 6
rect 1787 -19 1791 6
rect 1795 -19 1799 6
rect 1817 -19 1821 6
rect 1825 -19 1829 6
rect 1861 -19 1865 6
rect 1869 -19 1873 6
rect 1906 -19 1910 6
rect 1914 -19 1918 6
rect 1956 -21 1960 9
rect 1964 -21 1968 9
rect 1990 -21 1994 14
rect 1998 -21 2002 14
rect 2079 9 2083 21
rect 2087 9 2091 21
rect 2118 -7 2122 17
rect 2127 -7 2131 17
rect 2136 -7 2140 17
rect 2146 -13 2150 11
rect 2155 -13 2159 11
rect 2164 -13 2168 11
rect 2079 -46 2083 -34
rect 2087 -46 2091 -34
rect 2216 -15 2220 10
rect 2224 -15 2228 10
rect 2232 -15 2236 10
rect 2254 -15 2258 10
rect 2262 -15 2266 10
rect 2298 -15 2302 10
rect 2306 -15 2310 10
rect 2343 -15 2347 10
rect 2351 -15 2355 10
rect 2378 -15 2382 5
rect 2386 -15 2390 5
<< polysilicon >>
rect 1639 873 1641 876
rect 1647 873 1649 876
rect 1677 873 1679 876
rect 1721 873 1723 876
rect 1766 873 1768 876
rect 2179 874 2182 876
rect 2192 874 2210 876
rect 2230 874 2233 876
rect 1866 859 1868 862
rect 1876 859 1878 862
rect 1908 859 1910 862
rect 1639 841 1641 848
rect 1634 837 1641 841
rect 1635 826 1637 837
rect 1647 829 1649 848
rect 1677 840 1679 848
rect 1721 840 1723 848
rect 1671 838 1679 840
rect 1715 838 1723 840
rect 1671 826 1673 838
rect 1679 826 1681 835
rect 1715 826 1717 838
rect 1723 826 1725 835
rect 1766 826 1768 848
rect 1866 824 1868 847
rect 1876 824 1878 847
rect 1908 829 1910 847
rect 2217 836 2219 839
rect 2096 829 2098 836
rect 2103 829 2105 836
rect 2129 829 2131 836
rect 2156 829 2158 836
rect 2179 829 2181 836
rect 1635 813 1637 816
rect 1671 813 1673 816
rect 1679 813 1681 816
rect 1715 813 1717 816
rect 1723 813 1725 816
rect 1766 813 1768 816
rect 1908 819 1910 822
rect 1866 807 1868 811
rect 1876 807 1878 811
rect 2059 788 2061 791
rect 1855 770 1857 773
rect 1894 766 1896 769
rect 1904 766 1906 769
rect 2096 785 2098 788
rect 2103 785 2105 788
rect 2129 785 2131 789
rect 2156 785 2158 789
rect 2179 785 2181 789
rect 2217 781 2219 796
rect 2254 778 2256 781
rect 2300 777 2302 780
rect 2308 777 2310 780
rect 2338 777 2340 780
rect 2382 777 2384 780
rect 2427 777 2429 780
rect 1629 746 1631 749
rect 1637 746 1639 749
rect 1667 746 1669 749
rect 1711 746 1713 749
rect 1756 746 1758 749
rect 1855 744 1857 758
rect 1922 760 1924 763
rect 1932 760 1934 763
rect 1855 735 1857 738
rect 1894 733 1896 742
rect 1904 732 1906 742
rect 2059 750 2061 768
rect 2082 751 2084 758
rect 2106 751 2108 758
rect 2127 751 2129 758
rect 2144 751 2146 758
rect 2162 752 2164 759
rect 2201 757 2203 760
rect 2059 737 2061 740
rect 1629 714 1631 721
rect 1624 710 1631 714
rect 1625 699 1627 710
rect 1637 702 1639 721
rect 1667 713 1669 721
rect 1711 713 1713 721
rect 1661 711 1669 713
rect 1705 711 1713 713
rect 1661 699 1663 711
rect 1669 699 1671 708
rect 1705 699 1707 711
rect 1713 699 1715 708
rect 1756 699 1758 721
rect 1855 715 1857 718
rect 1855 689 1857 703
rect 1894 701 1896 728
rect 1904 701 1906 727
rect 1922 725 1924 736
rect 1922 701 1924 721
rect 1932 714 1934 736
rect 2254 753 2256 768
rect 2461 771 2463 774
rect 2300 745 2302 752
rect 2295 741 2302 745
rect 2201 719 2203 737
rect 2296 730 2298 741
rect 2308 733 2310 752
rect 2338 744 2340 752
rect 2382 744 2384 752
rect 2332 742 2340 744
rect 2376 742 2384 744
rect 2332 730 2334 742
rect 2340 730 2342 739
rect 2376 730 2378 742
rect 2384 730 2386 739
rect 2427 730 2429 752
rect 2461 733 2463 751
rect 2461 720 2463 723
rect 1932 701 1934 710
rect 2082 707 2084 711
rect 2106 707 2108 711
rect 2127 707 2129 711
rect 2144 707 2146 711
rect 2162 708 2164 712
rect 2296 717 2298 720
rect 2332 717 2334 720
rect 2340 717 2342 720
rect 2376 717 2378 720
rect 2384 717 2386 720
rect 2427 717 2429 720
rect 2201 706 2203 709
rect 1625 686 1627 689
rect 1661 686 1663 689
rect 1669 686 1671 689
rect 1705 686 1707 689
rect 1713 686 1715 689
rect 1756 686 1758 689
rect 1894 686 1896 689
rect 1904 686 1906 689
rect 1922 686 1924 689
rect 1932 686 1934 689
rect 2306 684 2308 687
rect 1855 680 1857 683
rect 2345 680 2347 683
rect 2355 680 2357 683
rect 2306 658 2308 672
rect 2373 674 2375 677
rect 2383 674 2385 677
rect 2306 649 2308 652
rect 2345 647 2347 656
rect 2355 646 2357 656
rect 2430 663 2432 666
rect 2438 663 2440 666
rect 2468 663 2470 666
rect 2512 663 2514 666
rect 2557 663 2559 666
rect 1640 639 1642 642
rect 1648 639 1650 642
rect 1678 639 1680 642
rect 1722 639 1724 642
rect 1767 639 1769 642
rect 2175 640 2178 642
rect 2188 640 2206 642
rect 2226 640 2229 642
rect 2306 629 2308 632
rect 1857 624 1859 627
rect 1867 624 1869 627
rect 1899 624 1901 627
rect 1640 607 1642 614
rect 1635 603 1642 607
rect 1636 592 1638 603
rect 1648 595 1650 614
rect 1678 606 1680 614
rect 1722 606 1724 614
rect 1672 604 1680 606
rect 1716 604 1724 606
rect 1672 592 1674 604
rect 1680 592 1682 601
rect 1716 592 1718 604
rect 1724 592 1726 601
rect 1767 592 1769 614
rect 2213 614 2215 617
rect 1857 589 1859 612
rect 1867 589 1869 612
rect 1899 594 1901 612
rect 2109 607 2111 614
rect 2116 607 2118 614
rect 2142 607 2144 614
rect 2169 607 2171 614
rect 1636 579 1638 582
rect 1672 579 1674 582
rect 1680 579 1682 582
rect 1716 579 1718 582
rect 1724 579 1726 582
rect 1767 579 1769 582
rect 1899 584 1901 587
rect 1857 572 1859 576
rect 1867 572 1869 576
rect 2072 565 2074 568
rect 2306 603 2308 617
rect 2345 615 2347 642
rect 2355 615 2357 641
rect 2373 639 2375 650
rect 2373 615 2375 635
rect 2383 628 2385 650
rect 2591 658 2593 661
rect 2430 631 2432 638
rect 2425 627 2432 631
rect 2383 615 2385 624
rect 2426 616 2428 627
rect 2438 619 2440 638
rect 2468 630 2470 638
rect 2512 630 2514 638
rect 2462 628 2470 630
rect 2506 628 2514 630
rect 2462 616 2464 628
rect 2470 616 2472 625
rect 2506 616 2508 628
rect 2514 616 2516 625
rect 2557 616 2559 638
rect 2591 620 2593 638
rect 2591 607 2593 610
rect 2426 603 2428 606
rect 2462 603 2464 606
rect 2470 603 2472 606
rect 2506 603 2508 606
rect 2514 603 2516 606
rect 2557 603 2559 606
rect 2345 600 2347 603
rect 2355 600 2357 603
rect 2373 600 2375 603
rect 2383 600 2385 603
rect 2306 594 2308 597
rect 2109 563 2111 566
rect 2116 563 2118 566
rect 2142 563 2144 567
rect 2169 563 2171 567
rect 2213 559 2215 574
rect 2250 556 2252 559
rect 1853 535 1855 538
rect 1892 531 1894 534
rect 1902 531 1904 534
rect 1645 514 1647 517
rect 1653 514 1655 517
rect 1683 514 1685 517
rect 1727 514 1729 517
rect 1772 514 1774 517
rect 1853 509 1855 523
rect 1920 525 1922 528
rect 1930 525 1932 528
rect 2072 527 2074 545
rect 2095 529 2097 536
rect 2119 529 2121 536
rect 2140 529 2142 536
rect 2157 529 2159 536
rect 2197 535 2199 538
rect 1853 500 1855 503
rect 1892 498 1894 507
rect 1902 497 1904 507
rect 2072 514 2074 517
rect 1645 482 1647 489
rect 1640 478 1647 482
rect 1641 467 1643 478
rect 1653 470 1655 489
rect 1683 481 1685 489
rect 1727 481 1729 489
rect 1677 479 1685 481
rect 1721 479 1729 481
rect 1677 467 1679 479
rect 1685 467 1687 476
rect 1721 467 1723 479
rect 1729 467 1731 476
rect 1772 467 1774 489
rect 1853 480 1855 483
rect 1641 454 1643 457
rect 1677 454 1679 457
rect 1685 454 1687 457
rect 1721 454 1723 457
rect 1729 454 1731 457
rect 1772 454 1774 457
rect 1853 454 1855 468
rect 1892 466 1894 493
rect 1902 466 1904 492
rect 1920 490 1922 501
rect 1920 466 1922 486
rect 1930 479 1932 501
rect 2250 531 2252 546
rect 2197 497 2199 515
rect 2095 485 2097 489
rect 2119 485 2121 489
rect 2140 485 2142 489
rect 2157 485 2159 489
rect 2305 492 2307 495
rect 2197 484 2199 487
rect 2344 488 2346 491
rect 2354 488 2356 491
rect 1930 466 1932 475
rect 2305 466 2307 480
rect 2372 482 2374 485
rect 2382 482 2384 485
rect 2305 457 2307 460
rect 2344 455 2346 464
rect 1892 451 1894 454
rect 1902 451 1904 454
rect 1920 451 1922 454
rect 1930 451 1932 454
rect 2354 454 2356 464
rect 2438 472 2440 475
rect 2446 472 2448 475
rect 2476 472 2478 475
rect 2520 472 2522 475
rect 2565 472 2567 475
rect 1853 445 1855 448
rect 2180 447 2183 449
rect 2193 447 2211 449
rect 2231 447 2234 449
rect 2305 437 2307 440
rect 1642 420 1644 423
rect 1650 420 1652 423
rect 1680 420 1682 423
rect 1724 420 1726 423
rect 1769 420 1771 423
rect 2218 420 2220 423
rect 2141 413 2143 420
rect 2148 413 2150 420
rect 2174 413 2176 420
rect 1865 405 1867 408
rect 1875 405 1877 408
rect 1907 405 1909 408
rect 1642 388 1644 395
rect 1637 384 1644 388
rect 1638 373 1640 384
rect 1650 376 1652 395
rect 1680 387 1682 395
rect 1724 387 1726 395
rect 1674 385 1682 387
rect 1718 385 1726 387
rect 1674 373 1676 385
rect 1682 373 1684 382
rect 1718 373 1720 385
rect 1726 373 1728 382
rect 1769 373 1771 395
rect 1865 370 1867 393
rect 1875 370 1877 393
rect 1907 375 1909 393
rect 1638 360 1640 363
rect 1674 360 1676 363
rect 1682 360 1684 363
rect 1718 360 1720 363
rect 1726 360 1728 363
rect 1769 360 1771 363
rect 2105 371 2107 374
rect 2305 411 2307 425
rect 2344 423 2346 450
rect 2354 423 2356 449
rect 2372 447 2374 458
rect 2372 423 2374 443
rect 2382 436 2384 458
rect 2598 467 2600 470
rect 2438 440 2440 447
rect 2433 436 2440 440
rect 2382 423 2384 432
rect 2434 425 2436 436
rect 2446 428 2448 447
rect 2476 439 2478 447
rect 2520 439 2522 447
rect 2470 437 2478 439
rect 2514 437 2522 439
rect 2470 425 2472 437
rect 2478 425 2480 434
rect 2514 425 2516 437
rect 2522 425 2524 434
rect 2565 425 2567 447
rect 2598 429 2600 447
rect 2598 416 2600 419
rect 2434 412 2436 415
rect 2470 412 2472 415
rect 2478 412 2480 415
rect 2514 412 2516 415
rect 2522 412 2524 415
rect 2565 412 2567 415
rect 2344 408 2346 411
rect 2354 408 2356 411
rect 2372 408 2374 411
rect 2382 408 2384 411
rect 2305 402 2307 405
rect 1907 365 1909 368
rect 1865 353 1867 357
rect 1875 353 1877 357
rect 2141 369 2143 372
rect 2148 369 2150 372
rect 2174 369 2176 373
rect 2218 365 2220 380
rect 2255 362 2257 365
rect 1850 332 1852 335
rect 2105 333 2107 351
rect 2127 335 2129 342
rect 2151 335 2153 342
rect 2172 335 2174 342
rect 2202 341 2204 344
rect 1889 328 1891 331
rect 1899 328 1901 331
rect 1653 306 1655 309
rect 1661 306 1663 309
rect 1691 306 1693 309
rect 1735 306 1737 309
rect 1780 306 1782 309
rect 1850 306 1852 320
rect 1917 322 1919 325
rect 1927 322 1929 325
rect 1850 297 1852 300
rect 1889 295 1891 304
rect 1899 294 1901 304
rect 2105 320 2107 323
rect 1653 274 1655 281
rect 1648 270 1655 274
rect 1649 259 1651 270
rect 1661 262 1663 281
rect 1691 273 1693 281
rect 1735 273 1737 281
rect 1685 271 1693 273
rect 1729 271 1737 273
rect 1685 259 1687 271
rect 1693 259 1695 268
rect 1729 259 1731 271
rect 1737 259 1739 268
rect 1780 259 1782 281
rect 1850 277 1852 280
rect 1850 251 1852 265
rect 1889 263 1891 290
rect 1899 263 1901 289
rect 1917 287 1919 298
rect 1917 263 1919 283
rect 1927 276 1929 298
rect 2255 337 2257 352
rect 2202 303 2204 321
rect 2127 291 2129 295
rect 2151 291 2153 295
rect 2172 291 2174 295
rect 2323 295 2325 298
rect 2202 290 2204 293
rect 2362 291 2364 294
rect 2372 291 2374 294
rect 1927 263 1929 272
rect 2323 269 2325 283
rect 2390 285 2392 288
rect 2400 285 2402 288
rect 2323 260 2325 263
rect 2362 258 2364 267
rect 2372 257 2374 267
rect 2459 278 2461 281
rect 2467 278 2469 281
rect 2497 278 2499 281
rect 2541 278 2543 281
rect 2586 278 2588 281
rect 1649 246 1651 249
rect 1685 246 1687 249
rect 1693 246 1695 249
rect 1729 246 1731 249
rect 1737 246 1739 249
rect 1780 246 1782 249
rect 1889 248 1891 251
rect 1899 248 1901 251
rect 1917 248 1919 251
rect 1927 248 1929 251
rect 1850 242 1852 245
rect 2323 240 2325 243
rect 1640 211 1642 214
rect 1648 211 1650 214
rect 1678 211 1680 214
rect 1722 211 1724 214
rect 1767 211 1769 214
rect 1863 213 1865 216
rect 1873 213 1875 216
rect 1905 213 1907 216
rect 2323 214 2325 228
rect 2362 226 2364 253
rect 2372 226 2374 252
rect 2390 250 2392 261
rect 2390 226 2392 246
rect 2400 239 2402 261
rect 2621 273 2623 276
rect 2459 246 2461 253
rect 2454 242 2461 246
rect 2400 226 2402 235
rect 2455 231 2457 242
rect 2467 234 2469 253
rect 2497 245 2499 253
rect 2541 245 2543 253
rect 2491 243 2499 245
rect 2535 243 2543 245
rect 2491 231 2493 243
rect 2499 231 2501 240
rect 2535 231 2537 243
rect 2543 231 2545 240
rect 2586 231 2588 253
rect 2621 235 2623 253
rect 2621 222 2623 225
rect 2455 218 2457 221
rect 2491 218 2493 221
rect 2499 218 2501 221
rect 2535 218 2537 221
rect 2543 218 2545 221
rect 2586 218 2588 221
rect 2182 209 2185 211
rect 2195 209 2213 211
rect 2233 209 2236 211
rect 2362 211 2364 214
rect 2372 211 2374 214
rect 2390 211 2392 214
rect 2400 211 2402 214
rect 2323 205 2325 208
rect 1640 179 1642 186
rect 1635 175 1642 179
rect 1636 164 1638 175
rect 1648 167 1650 186
rect 1678 178 1680 186
rect 1722 178 1724 186
rect 1672 176 1680 178
rect 1716 176 1724 178
rect 1672 164 1674 176
rect 1680 164 1682 173
rect 1716 164 1718 176
rect 1724 164 1726 173
rect 1767 164 1769 186
rect 1863 178 1865 201
rect 1873 178 1875 201
rect 1905 183 1907 201
rect 2220 182 2222 185
rect 1905 173 1907 176
rect 2162 175 2164 182
rect 2169 175 2171 182
rect 1863 161 1865 165
rect 1873 161 1875 165
rect 1636 151 1638 154
rect 1672 151 1674 154
rect 1680 151 1682 154
rect 1716 151 1718 154
rect 1724 151 1726 154
rect 1767 151 1769 154
rect 1849 136 1851 139
rect 1888 132 1890 135
rect 1898 132 1900 135
rect 2124 134 2126 137
rect 1645 113 1647 116
rect 1653 113 1655 116
rect 1683 113 1685 116
rect 1727 113 1729 116
rect 1772 113 1774 116
rect 1849 110 1851 124
rect 1916 126 1918 129
rect 1926 126 1928 129
rect 1849 101 1851 104
rect 1888 99 1890 108
rect 1898 98 1900 108
rect 2162 131 2164 134
rect 2169 131 2171 134
rect 2220 127 2222 142
rect 2257 124 2259 127
rect 1645 81 1647 88
rect 1640 77 1647 81
rect 1641 66 1643 77
rect 1653 69 1655 88
rect 1683 80 1685 88
rect 1727 80 1729 88
rect 1677 78 1685 80
rect 1721 78 1729 80
rect 1677 66 1679 78
rect 1685 66 1687 75
rect 1721 66 1723 78
rect 1729 66 1731 75
rect 1772 66 1774 88
rect 1849 81 1851 84
rect 1641 53 1643 56
rect 1677 53 1679 56
rect 1685 53 1687 56
rect 1721 53 1723 56
rect 1729 53 1731 56
rect 1772 53 1774 56
rect 1849 55 1851 69
rect 1888 67 1890 94
rect 1898 67 1900 93
rect 1916 91 1918 102
rect 1916 67 1918 87
rect 1926 80 1928 102
rect 2124 96 2126 114
rect 2148 97 2150 104
rect 2172 97 2174 104
rect 2204 103 2206 106
rect 2124 83 2126 86
rect 1926 67 1928 76
rect 2257 99 2259 114
rect 2204 65 2206 83
rect 1888 52 1890 55
rect 1898 52 1900 55
rect 1916 52 1918 55
rect 1926 52 1928 55
rect 2148 53 2150 57
rect 2172 53 2174 57
rect 2204 52 2206 55
rect 1849 46 1851 49
rect 2084 21 2086 24
rect 1995 14 1997 17
rect 1961 9 1963 12
rect 1784 6 1786 9
rect 1792 6 1794 9
rect 1822 6 1824 9
rect 1866 6 1868 9
rect 1911 6 1913 9
rect 1784 -26 1786 -19
rect 1779 -30 1786 -26
rect 1780 -41 1782 -30
rect 1792 -38 1794 -19
rect 1822 -27 1824 -19
rect 1866 -27 1868 -19
rect 1816 -29 1824 -27
rect 1860 -29 1868 -27
rect 1816 -41 1818 -29
rect 1824 -41 1826 -32
rect 1860 -41 1862 -29
rect 1868 -41 1870 -32
rect 1911 -41 1913 -19
rect 2123 17 2125 20
rect 2133 17 2135 20
rect 2084 -5 2086 9
rect 2151 11 2153 14
rect 2161 11 2163 14
rect 2084 -14 2086 -11
rect 2123 -16 2125 -7
rect 2133 -17 2135 -7
rect 2221 10 2223 13
rect 2229 10 2231 13
rect 2259 10 2261 13
rect 2303 10 2305 13
rect 2348 10 2350 13
rect 1961 -39 1963 -21
rect 1995 -39 1997 -21
rect 2084 -34 2086 -31
rect 1780 -54 1782 -51
rect 1816 -54 1818 -51
rect 1824 -54 1826 -51
rect 1860 -54 1862 -51
rect 1868 -54 1870 -51
rect 1911 -54 1913 -51
rect 1961 -58 1963 -55
rect 1995 -61 1997 -58
rect 2084 -60 2086 -46
rect 2123 -48 2125 -21
rect 2133 -48 2135 -22
rect 2151 -24 2153 -13
rect 2151 -48 2153 -28
rect 2161 -35 2163 -13
rect 2383 5 2385 8
rect 2221 -22 2223 -15
rect 2216 -26 2223 -22
rect 2217 -37 2219 -26
rect 2229 -34 2231 -15
rect 2259 -23 2261 -15
rect 2303 -23 2305 -15
rect 2253 -25 2261 -23
rect 2297 -25 2305 -23
rect 2253 -37 2255 -25
rect 2261 -37 2263 -28
rect 2297 -37 2299 -25
rect 2305 -37 2307 -28
rect 2348 -37 2350 -15
rect 2383 -33 2385 -15
rect 2161 -48 2163 -39
rect 2383 -46 2385 -43
rect 2217 -50 2219 -47
rect 2253 -50 2255 -47
rect 2261 -50 2263 -47
rect 2297 -50 2299 -47
rect 2305 -50 2307 -47
rect 2348 -50 2350 -47
rect 2123 -63 2125 -60
rect 2133 -63 2135 -60
rect 2151 -63 2153 -60
rect 2161 -63 2163 -60
rect 2084 -69 2086 -66
<< polycontact >>
rect 2196 876 2200 880
rect 1630 837 1634 841
rect 1643 829 1647 833
rect 1654 837 1658 841
rect 1666 829 1671 834
rect 1681 829 1685 833
rect 1710 829 1715 834
rect 1762 834 1766 839
rect 1725 829 1729 833
rect 1862 834 1866 838
rect 1872 827 1876 831
rect 1904 833 1908 837
rect 2092 832 2096 836
rect 2105 832 2109 836
rect 2125 832 2129 836
rect 2152 832 2156 836
rect 2175 832 2179 836
rect 2213 781 2217 785
rect 1851 747 1855 751
rect 2055 754 2059 758
rect 2078 754 2082 758
rect 2102 754 2106 758
rect 2123 754 2127 758
rect 2140 754 2144 758
rect 2158 755 2162 759
rect 1620 710 1624 714
rect 1633 702 1637 706
rect 1644 710 1648 714
rect 1656 702 1661 707
rect 1671 702 1675 706
rect 1700 702 1705 707
rect 1752 707 1756 712
rect 1715 702 1719 706
rect 1851 692 1855 696
rect 1920 721 1924 725
rect 1931 710 1935 714
rect 2250 753 2254 757
rect 2291 741 2295 745
rect 2197 723 2201 727
rect 2304 733 2308 737
rect 2315 741 2319 745
rect 2327 733 2332 738
rect 2342 733 2346 737
rect 2371 733 2376 738
rect 2423 738 2427 743
rect 2386 733 2390 737
rect 2457 737 2461 741
rect 2302 661 2306 665
rect 2192 642 2196 646
rect 1631 603 1635 607
rect 1644 595 1648 599
rect 1655 603 1659 607
rect 1667 595 1672 600
rect 1682 595 1686 599
rect 1711 595 1716 600
rect 1763 600 1767 605
rect 1726 595 1730 599
rect 1853 599 1857 603
rect 1863 592 1867 596
rect 1895 598 1899 602
rect 2105 610 2109 614
rect 2118 610 2122 614
rect 2138 610 2142 614
rect 2165 610 2169 614
rect 2302 606 2306 610
rect 2371 635 2375 639
rect 2382 624 2386 628
rect 2421 627 2425 631
rect 2434 619 2438 623
rect 2445 627 2449 631
rect 2457 619 2462 624
rect 2472 619 2476 623
rect 2501 619 2506 624
rect 2553 624 2557 629
rect 2516 619 2520 623
rect 2587 624 2591 628
rect 2209 559 2213 563
rect 2068 531 2072 535
rect 1849 512 1853 516
rect 2091 532 2095 536
rect 2115 532 2119 536
rect 2136 532 2140 536
rect 2153 532 2157 536
rect 1636 478 1640 482
rect 1649 470 1653 474
rect 1660 478 1664 482
rect 1672 470 1677 475
rect 1687 470 1691 474
rect 1716 470 1721 475
rect 1768 475 1772 480
rect 1731 470 1735 474
rect 1849 457 1853 461
rect 1918 486 1922 490
rect 2246 531 2250 535
rect 2193 501 2197 505
rect 1929 475 1933 479
rect 2301 469 2305 473
rect 2197 449 2201 453
rect 2137 416 2141 420
rect 2150 416 2154 420
rect 2170 416 2174 420
rect 1633 384 1637 388
rect 1646 376 1650 380
rect 1657 384 1661 388
rect 1669 376 1674 381
rect 1684 376 1688 380
rect 1713 376 1718 381
rect 1765 381 1769 386
rect 1728 376 1732 380
rect 1861 380 1865 384
rect 1871 373 1875 377
rect 1903 379 1907 383
rect 2301 414 2305 418
rect 2370 443 2374 447
rect 2429 436 2433 440
rect 2381 432 2385 436
rect 2442 428 2446 432
rect 2453 436 2457 440
rect 2465 428 2470 433
rect 2480 428 2484 432
rect 2509 428 2514 433
rect 2561 433 2565 438
rect 2524 428 2528 432
rect 2594 433 2598 437
rect 2214 365 2218 369
rect 2101 337 2105 341
rect 2123 338 2127 342
rect 2147 338 2151 342
rect 2168 338 2172 342
rect 1846 309 1850 313
rect 1644 270 1648 274
rect 1657 262 1661 266
rect 1668 270 1672 274
rect 1680 262 1685 267
rect 1695 262 1699 266
rect 1724 262 1729 267
rect 1776 267 1780 272
rect 1739 262 1743 266
rect 1846 254 1850 258
rect 1915 283 1919 287
rect 2251 337 2255 341
rect 2198 307 2202 311
rect 1926 272 1930 276
rect 2319 272 2323 276
rect 2319 217 2323 221
rect 2199 211 2203 215
rect 2388 246 2392 250
rect 2450 242 2454 246
rect 2399 235 2403 239
rect 2463 234 2467 238
rect 2474 242 2478 246
rect 2486 234 2491 239
rect 2501 234 2505 238
rect 2530 234 2535 239
rect 2582 239 2586 244
rect 2545 234 2549 238
rect 2617 239 2621 243
rect 1859 188 1863 192
rect 1631 175 1635 179
rect 1644 167 1648 171
rect 1655 175 1659 179
rect 1667 167 1672 172
rect 1682 167 1686 171
rect 1711 167 1716 172
rect 1763 172 1767 177
rect 1726 167 1730 171
rect 1869 181 1873 185
rect 1901 187 1905 191
rect 2158 178 2162 182
rect 2171 178 2175 182
rect 1845 113 1849 117
rect 2216 127 2220 131
rect 1636 77 1640 81
rect 1649 69 1653 73
rect 1660 77 1664 81
rect 1672 69 1677 74
rect 1687 69 1691 73
rect 1716 69 1721 74
rect 1768 74 1772 79
rect 1731 69 1735 73
rect 1845 58 1849 62
rect 1914 87 1918 91
rect 2120 100 2124 104
rect 2144 100 2148 104
rect 2168 100 2172 104
rect 1925 76 1929 80
rect 2253 99 2257 103
rect 2200 69 2204 73
rect 1775 -30 1779 -26
rect 1788 -38 1792 -34
rect 1799 -30 1803 -26
rect 1811 -38 1816 -33
rect 1826 -38 1830 -34
rect 1855 -38 1860 -33
rect 1907 -33 1911 -28
rect 1870 -38 1874 -34
rect 2080 -2 2084 2
rect 1957 -35 1961 -31
rect 1991 -35 1995 -31
rect 2080 -57 2084 -53
rect 2149 -28 2153 -24
rect 2212 -26 2216 -22
rect 2160 -39 2164 -35
rect 2225 -34 2229 -30
rect 2236 -26 2240 -22
rect 2248 -34 2253 -29
rect 2263 -34 2267 -30
rect 2292 -34 2297 -29
rect 2344 -29 2348 -24
rect 2307 -34 2311 -30
rect 2379 -29 2383 -25
<< metal1 >>
rect 1628 879 1781 883
rect 1634 873 1638 879
rect 1672 873 1676 879
rect 1716 873 1720 879
rect 1761 873 1765 879
rect 1684 848 1697 873
rect 1728 848 1741 873
rect 1966 870 1969 903
rect 1853 865 1924 868
rect 1623 837 1630 841
rect 1634 829 1643 833
rect 1650 826 1654 848
rect 1658 837 1659 841
rect 1694 839 1697 848
rect 1738 839 1741 848
rect 1694 834 1706 839
rect 1738 834 1762 839
rect 1769 838 1773 848
rect 1861 859 1865 865
rect 1879 859 1883 865
rect 1903 859 1906 865
rect 1870 844 1873 847
rect 1870 841 1883 844
rect 1769 834 1862 838
rect 1880 837 1883 841
rect 1912 837 1915 847
rect 1658 832 1666 834
rect 1663 829 1666 832
rect 1685 829 1686 833
rect 1694 826 1697 834
rect 1702 829 1710 834
rect 1729 829 1730 833
rect 1738 826 1741 834
rect 1769 833 1850 834
rect 1880 833 1904 837
rect 1912 834 1961 837
rect 1769 826 1773 833
rect 1642 816 1654 826
rect 1686 816 1697 826
rect 1730 816 1741 826
rect 1630 811 1634 816
rect 1666 811 1670 816
rect 1710 811 1714 816
rect 1761 811 1765 816
rect 1629 807 1773 811
rect 1618 752 1771 756
rect 1624 746 1628 752
rect 1662 746 1666 752
rect 1706 746 1710 752
rect 1751 746 1755 752
rect 1798 751 1803 833
rect 1857 830 1872 831
rect 1815 827 1872 830
rect 1815 760 1818 827
rect 1880 824 1883 833
rect 1912 829 1915 834
rect 1861 805 1864 811
rect 1903 805 1906 822
rect 1853 802 1906 805
rect 1849 776 1877 779
rect 1850 770 1853 776
rect 1874 775 1877 776
rect 1874 772 1945 775
rect 1798 749 1833 751
rect 1798 746 1836 749
rect 1674 721 1687 746
rect 1718 721 1731 746
rect 1841 747 1851 750
rect 1859 750 1862 758
rect 1889 766 1892 772
rect 1908 766 1911 772
rect 1859 747 1880 750
rect 1859 744 1862 747
rect 1613 710 1620 714
rect 1624 702 1633 706
rect 1640 699 1644 721
rect 1648 710 1649 714
rect 1684 712 1687 721
rect 1728 712 1731 721
rect 1684 707 1696 712
rect 1728 707 1752 712
rect 1759 711 1763 721
rect 1648 705 1656 707
rect 1653 702 1656 705
rect 1675 702 1676 706
rect 1684 699 1687 707
rect 1692 702 1700 707
rect 1719 702 1720 706
rect 1728 699 1731 707
rect 1759 706 1772 711
rect 1759 699 1763 706
rect 1632 689 1644 699
rect 1676 689 1687 699
rect 1720 689 1731 699
rect 1768 695 1771 706
rect 1815 695 1818 738
rect 1850 734 1853 738
rect 1844 732 1868 734
rect 1844 731 1862 732
rect 1867 731 1868 732
rect 1877 724 1880 747
rect 1918 766 1938 769
rect 1918 760 1921 766
rect 1935 760 1938 766
rect 1899 739 1902 742
rect 1899 736 1917 739
rect 1927 729 1930 736
rect 1927 726 1944 729
rect 1849 723 1868 724
rect 1844 721 1868 723
rect 1877 721 1920 724
rect 1850 715 1853 721
rect 1941 716 1944 726
rect 1906 710 1931 713
rect 1906 708 1909 710
rect 1768 692 1836 695
rect 1841 692 1851 695
rect 1859 695 1862 703
rect 1871 705 1909 708
rect 1941 707 1944 711
rect 1871 695 1874 705
rect 1912 704 1944 707
rect 1912 701 1915 704
rect 1859 692 1874 695
rect 1859 689 1862 692
rect 1620 684 1624 689
rect 1656 684 1660 689
rect 1700 684 1704 689
rect 1751 684 1755 689
rect 1619 680 1763 684
rect 1911 698 1917 701
rect 1850 679 1853 683
rect 1871 682 1876 685
rect 1889 685 1892 689
rect 1936 685 1939 689
rect 1881 682 1945 685
rect 1871 679 1874 682
rect 1844 676 1874 679
rect 1958 671 1961 834
rect 1966 717 1969 865
rect 1982 861 1986 904
rect 1966 660 1969 711
rect 1974 680 1977 805
rect 1629 645 1782 649
rect 1635 639 1639 645
rect 1673 639 1677 645
rect 1717 639 1721 645
rect 1762 639 1766 645
rect 1685 614 1698 639
rect 1729 614 1742 639
rect 1844 630 1915 633
rect 1624 603 1631 607
rect 1635 595 1644 599
rect 1651 592 1655 614
rect 1659 603 1660 607
rect 1695 605 1698 614
rect 1739 605 1742 614
rect 1695 600 1707 605
rect 1739 600 1763 605
rect 1770 604 1774 614
rect 1852 624 1856 630
rect 1870 624 1874 630
rect 1894 624 1897 630
rect 1861 609 1864 612
rect 1861 606 1874 609
rect 1770 603 1783 604
rect 1659 598 1667 600
rect 1664 595 1667 598
rect 1686 595 1687 599
rect 1695 592 1698 600
rect 1703 595 1711 600
rect 1730 595 1731 599
rect 1739 592 1742 600
rect 1770 599 1853 603
rect 1871 602 1874 606
rect 1903 602 1906 612
rect 1974 602 1977 675
rect 1982 641 1986 856
rect 1998 851 2002 903
rect 1991 689 1994 806
rect 1770 592 1774 599
rect 1643 582 1655 592
rect 1687 582 1698 592
rect 1731 582 1742 592
rect 1631 577 1635 582
rect 1667 577 1671 582
rect 1711 577 1715 582
rect 1762 577 1766 582
rect 1630 573 1774 577
rect 1634 520 1787 524
rect 1640 514 1644 520
rect 1678 514 1682 520
rect 1722 514 1726 520
rect 1767 514 1771 520
rect 1690 489 1703 514
rect 1734 489 1747 514
rect 1796 513 1800 599
rect 1871 598 1895 602
rect 1903 599 1977 602
rect 1819 592 1863 596
rect 1819 526 1823 592
rect 1871 589 1874 598
rect 1903 594 1906 599
rect 1852 570 1855 576
rect 1894 570 1897 587
rect 1844 567 1897 570
rect 1847 541 1875 544
rect 1848 535 1851 541
rect 1872 540 1875 541
rect 1872 537 1943 540
rect 1819 524 1824 526
rect 1812 514 1830 515
rect 1812 513 1834 514
rect 1796 511 1834 513
rect 1796 510 1830 511
rect 1839 512 1849 515
rect 1857 515 1860 523
rect 1887 531 1890 537
rect 1906 531 1909 537
rect 1857 512 1878 515
rect 1796 509 1814 510
rect 1857 509 1860 512
rect 1629 478 1636 482
rect 1640 470 1649 474
rect 1656 467 1660 489
rect 1664 478 1665 482
rect 1700 480 1703 489
rect 1744 480 1747 489
rect 1700 475 1712 480
rect 1744 475 1768 480
rect 1775 479 1779 489
rect 1819 479 1824 502
rect 1848 499 1851 503
rect 1842 497 1866 499
rect 1842 496 1860 497
rect 1865 496 1866 497
rect 1875 489 1878 512
rect 1916 531 1936 534
rect 1916 525 1919 531
rect 1933 525 1936 531
rect 1897 504 1900 507
rect 1897 501 1915 504
rect 1925 494 1928 501
rect 1974 494 1977 599
rect 1925 491 1942 494
rect 1847 488 1866 489
rect 1842 486 1866 488
rect 1875 486 1918 489
rect 1664 473 1672 475
rect 1669 470 1672 473
rect 1691 470 1692 474
rect 1700 467 1703 475
rect 1708 470 1716 475
rect 1735 470 1736 474
rect 1744 467 1747 475
rect 1775 474 1824 479
rect 1848 480 1851 486
rect 1939 480 1942 491
rect 1974 483 1977 489
rect 1982 484 1986 636
rect 1991 554 1994 684
rect 1998 632 2002 845
rect 2018 842 2022 901
rect 2007 698 2010 805
rect 2010 693 2011 698
rect 1981 480 1986 484
rect 1775 467 1779 474
rect 1648 457 1660 467
rect 1692 457 1703 467
rect 1736 457 1747 467
rect 1817 461 1822 474
rect 1904 475 1929 478
rect 1939 476 1987 480
rect 1904 473 1907 475
rect 1636 452 1640 457
rect 1672 452 1676 457
rect 1716 452 1720 457
rect 1767 452 1771 457
rect 1817 456 1834 461
rect 1839 457 1849 460
rect 1857 460 1860 468
rect 1869 470 1907 473
rect 1939 472 1942 476
rect 1869 460 1872 470
rect 1910 469 1942 472
rect 1981 472 1985 476
rect 1910 466 1913 469
rect 1857 457 1872 460
rect 1857 454 1860 457
rect 1635 448 1779 452
rect 1909 463 1915 466
rect 1981 465 1985 467
rect 1848 444 1851 448
rect 1869 447 1874 450
rect 1887 450 1890 454
rect 1934 450 1937 454
rect 1879 447 1943 450
rect 1869 444 1872 447
rect 1842 441 1872 444
rect 1631 426 1784 430
rect 1637 420 1641 426
rect 1675 420 1679 426
rect 1719 420 1723 426
rect 1764 420 1768 426
rect 1687 395 1700 420
rect 1731 395 1744 420
rect 1852 411 1923 414
rect 1626 384 1633 388
rect 1637 376 1646 380
rect 1653 373 1657 395
rect 1661 384 1662 388
rect 1697 386 1700 395
rect 1741 386 1744 395
rect 1697 381 1709 386
rect 1741 381 1765 386
rect 1772 385 1776 395
rect 1860 405 1864 411
rect 1878 405 1882 411
rect 1902 405 1905 411
rect 1991 396 1994 549
rect 1998 439 2002 627
rect 2007 544 2010 693
rect 2018 622 2022 837
rect 2033 835 2038 902
rect 2171 881 2174 888
rect 2171 878 2182 881
rect 2196 880 2200 888
rect 2236 881 2239 888
rect 2230 878 2239 881
rect 2192 869 2210 872
rect 2111 836 2115 837
rect 2089 835 2092 836
rect 2033 832 2092 835
rect 2109 832 2115 836
rect 2122 832 2125 845
rect 2147 836 2150 856
rect 2169 836 2173 865
rect 2197 860 2200 869
rect 2236 860 2239 878
rect 2147 832 2152 836
rect 2169 832 2175 836
rect 2182 835 2186 836
rect 1990 393 1995 396
rect 1869 390 1872 393
rect 1869 387 1882 390
rect 1772 384 1852 385
rect 1661 379 1669 381
rect 1666 376 1669 379
rect 1688 376 1689 380
rect 1697 373 1700 381
rect 1705 376 1713 381
rect 1732 376 1733 380
rect 1741 373 1744 381
rect 1772 380 1861 384
rect 1879 383 1882 387
rect 1911 383 1914 393
rect 1991 383 1994 393
rect 1772 373 1776 380
rect 1645 363 1657 373
rect 1689 363 1700 373
rect 1733 363 1744 373
rect 1633 358 1637 363
rect 1669 358 1673 363
rect 1713 358 1717 363
rect 1764 358 1768 363
rect 1632 354 1776 358
rect 1642 312 1795 316
rect 1648 306 1652 312
rect 1686 306 1690 312
rect 1730 306 1734 312
rect 1775 306 1779 312
rect 1798 310 1803 380
rect 1879 379 1903 383
rect 1911 380 1994 383
rect 1818 373 1871 377
rect 1818 321 1822 373
rect 1879 370 1882 379
rect 1911 375 1914 380
rect 1860 351 1863 357
rect 1902 351 1905 368
rect 1991 358 1994 380
rect 1852 348 1905 351
rect 1844 338 1872 341
rect 1845 332 1848 338
rect 1869 337 1872 338
rect 1869 334 1940 337
rect 1818 320 1821 321
rect 1809 310 1831 311
rect 1798 308 1831 310
rect 1798 306 1827 308
rect 1836 309 1846 312
rect 1854 312 1857 320
rect 1884 328 1887 334
rect 1903 328 1906 334
rect 1854 309 1875 312
rect 1854 306 1857 309
rect 1698 281 1711 306
rect 1742 281 1755 306
rect 1798 305 1813 306
rect 1637 270 1644 274
rect 1648 262 1657 266
rect 1664 259 1668 281
rect 1672 270 1673 274
rect 1708 272 1711 281
rect 1752 272 1755 281
rect 1708 267 1720 272
rect 1752 267 1776 272
rect 1783 271 1787 281
rect 1816 271 1821 298
rect 1845 296 1848 300
rect 1839 294 1863 296
rect 1839 293 1857 294
rect 1862 293 1863 294
rect 1872 286 1875 309
rect 1913 328 1933 331
rect 1913 322 1916 328
rect 1930 322 1933 328
rect 1894 301 1897 304
rect 1894 298 1912 301
rect 1922 291 1925 298
rect 1991 296 1994 353
rect 1998 293 2002 434
rect 2007 350 2010 539
rect 2018 429 2022 617
rect 1922 288 1939 291
rect 1844 285 1863 286
rect 1839 283 1863 285
rect 1872 283 1915 286
rect 1672 265 1680 267
rect 1677 262 1680 265
rect 1699 262 1700 266
rect 1708 259 1711 267
rect 1716 262 1724 267
rect 1743 262 1744 266
rect 1752 259 1755 267
rect 1783 266 1821 271
rect 1783 259 1787 266
rect 1656 249 1668 259
rect 1700 249 1711 259
rect 1744 249 1755 259
rect 1818 257 1821 266
rect 1845 277 1848 283
rect 1936 277 1939 288
rect 1998 277 2001 293
rect 1901 272 1926 275
rect 1936 274 2001 277
rect 1901 270 1904 272
rect 1818 254 1831 257
rect 1836 254 1846 257
rect 1854 257 1857 265
rect 1866 267 1904 270
rect 1936 269 1939 274
rect 1866 257 1869 267
rect 1907 266 1939 269
rect 1998 266 2001 274
rect 1907 263 1910 266
rect 1854 254 1869 257
rect 1854 251 1857 254
rect 1644 244 1648 249
rect 1680 244 1684 249
rect 1724 244 1728 249
rect 1775 244 1779 249
rect 1906 260 1912 263
rect 1643 240 1787 244
rect 1845 241 1848 245
rect 1866 244 1871 247
rect 1884 247 1887 251
rect 1931 247 1934 251
rect 1876 244 1940 247
rect 1866 241 1869 244
rect 1839 238 1869 241
rect 1629 217 1782 221
rect 1850 219 1921 222
rect 1635 211 1639 217
rect 1673 211 1677 217
rect 1717 211 1721 217
rect 1762 211 1766 217
rect 1858 213 1862 219
rect 1876 213 1880 219
rect 1685 186 1698 211
rect 1729 186 1742 211
rect 1900 213 1903 219
rect 1998 201 2001 261
rect 1867 198 1870 201
rect 1867 195 1880 198
rect 1826 192 1852 193
rect 1624 175 1631 179
rect 1635 167 1644 171
rect 1651 164 1655 186
rect 1659 175 1660 179
rect 1695 177 1698 186
rect 1739 177 1742 186
rect 1695 172 1707 177
rect 1739 172 1763 177
rect 1770 176 1774 186
rect 1800 188 1859 192
rect 1877 191 1880 195
rect 1909 191 1912 201
rect 2007 191 2010 345
rect 1800 187 1826 188
rect 1877 187 1901 191
rect 1909 188 2010 191
rect 2018 191 2022 424
rect 2033 613 2038 832
rect 2182 831 2193 835
rect 2182 829 2186 831
rect 2047 794 2075 797
rect 2054 788 2057 794
rect 2091 779 2095 788
rect 2106 787 2111 788
rect 2124 787 2128 789
rect 2106 782 2128 787
rect 2132 787 2136 789
rect 2151 787 2155 789
rect 2132 782 2155 787
rect 2159 787 2163 789
rect 2174 787 2178 789
rect 2159 782 2178 787
rect 2086 775 2104 779
rect 2063 758 2066 768
rect 2047 754 2055 758
rect 2063 755 2078 758
rect 2063 750 2066 755
rect 2075 754 2078 755
rect 2085 751 2089 760
rect 2054 732 2057 740
rect 2047 729 2057 732
rect 2077 706 2081 711
rect 2092 706 2096 775
rect 2099 754 2102 764
rect 2109 751 2113 782
rect 2137 778 2141 782
rect 2164 779 2168 782
rect 2189 780 2193 831
rect 2196 785 2200 860
rect 2205 842 2233 845
rect 2212 836 2215 842
rect 2196 781 2213 785
rect 2221 784 2224 796
rect 2236 791 2277 794
rect 2236 784 2239 791
rect 2242 784 2270 787
rect 2221 781 2239 784
rect 2130 774 2141 778
rect 2147 775 2168 779
rect 2181 778 2193 780
rect 2225 778 2229 781
rect 2181 776 2229 778
rect 2120 754 2123 764
rect 2130 751 2134 774
rect 2137 754 2140 762
rect 2147 751 2151 775
rect 2155 769 2160 770
rect 2155 755 2158 764
rect 2181 759 2185 776
rect 2189 774 2229 776
rect 2249 778 2252 784
rect 2189 763 2217 766
rect 2165 755 2185 759
rect 2165 752 2169 755
rect 2181 727 2185 755
rect 2196 757 2199 763
rect 2220 754 2250 757
rect 2220 745 2223 754
rect 2242 753 2250 754
rect 2258 756 2261 768
rect 2274 756 2277 791
rect 2289 783 2442 787
rect 2258 753 2277 756
rect 2295 777 2299 783
rect 2333 777 2337 783
rect 2377 777 2381 783
rect 2422 777 2426 783
rect 2449 777 2477 780
rect 2345 752 2358 777
rect 2389 752 2402 777
rect 2219 741 2291 745
rect 2205 727 2208 737
rect 2220 727 2223 741
rect 2295 733 2304 737
rect 2311 730 2315 752
rect 2319 741 2320 745
rect 2355 743 2358 752
rect 2399 743 2402 752
rect 2355 738 2367 743
rect 2399 738 2423 743
rect 2430 742 2434 752
rect 2456 771 2459 777
rect 2430 741 2443 742
rect 2465 741 2468 751
rect 2319 736 2327 738
rect 2324 733 2327 736
rect 2346 733 2347 737
rect 2355 730 2358 738
rect 2363 733 2371 738
rect 2390 733 2391 737
rect 2399 730 2402 738
rect 2430 737 2457 741
rect 2465 738 2477 741
rect 2430 730 2434 737
rect 2465 733 2468 738
rect 2181 723 2197 727
rect 2205 724 2223 727
rect 2205 719 2208 724
rect 2101 706 2105 711
rect 2122 706 2126 711
rect 2139 706 2143 711
rect 2157 706 2161 712
rect 2077 703 2161 706
rect 2303 720 2315 730
rect 2347 720 2358 730
rect 2391 720 2402 730
rect 2291 715 2295 720
rect 2327 715 2331 720
rect 2371 715 2375 720
rect 2422 715 2426 720
rect 2456 715 2459 723
rect 2290 711 2434 715
rect 2449 712 2459 715
rect 2196 701 2199 709
rect 2185 698 2199 701
rect 2300 690 2328 693
rect 2301 684 2304 690
rect 2325 689 2328 690
rect 2325 686 2396 689
rect 2274 662 2287 663
rect 2279 660 2287 662
rect 2292 661 2302 664
rect 2310 664 2313 672
rect 2340 680 2343 686
rect 2359 680 2362 686
rect 2310 661 2331 664
rect 2310 658 2313 661
rect 2167 647 2170 654
rect 2167 644 2178 647
rect 2192 646 2196 654
rect 2232 647 2235 654
rect 2301 648 2304 652
rect 2226 644 2235 647
rect 2295 646 2319 648
rect 2295 645 2313 646
rect 2157 639 2158 641
rect 2157 636 2165 639
rect 2139 627 2140 632
rect 2124 614 2128 617
rect 2102 613 2105 614
rect 2033 610 2105 613
rect 2122 610 2128 614
rect 2135 610 2138 627
rect 2162 610 2165 636
rect 2188 635 2206 638
rect 2193 626 2196 635
rect 2232 626 2235 644
rect 2318 645 2319 646
rect 2328 638 2331 661
rect 2369 680 2389 683
rect 2369 674 2372 680
rect 2386 674 2389 680
rect 2350 653 2353 656
rect 2350 650 2368 653
rect 2419 669 2572 673
rect 2425 663 2429 669
rect 2463 663 2467 669
rect 2507 663 2511 669
rect 2552 663 2556 669
rect 2579 664 2607 667
rect 2378 643 2381 650
rect 2378 640 2395 643
rect 2300 637 2319 638
rect 2295 635 2319 637
rect 2328 635 2371 638
rect 2301 629 2304 635
rect 2392 631 2395 640
rect 2475 638 2488 663
rect 2519 638 2532 663
rect 2586 658 2589 664
rect 2033 419 2038 610
rect 2060 571 2088 574
rect 2067 565 2070 571
rect 2104 557 2108 566
rect 2119 565 2124 566
rect 2137 565 2141 567
rect 2119 560 2141 565
rect 2145 565 2149 567
rect 2164 565 2168 567
rect 2145 560 2168 565
rect 2172 565 2176 567
rect 2172 560 2181 565
rect 2103 553 2110 557
rect 2076 535 2079 545
rect 2088 535 2091 536
rect 2060 531 2068 535
rect 2076 532 2091 535
rect 2076 527 2079 532
rect 2098 529 2102 538
rect 2067 509 2070 517
rect 2060 506 2070 509
rect 2090 484 2094 489
rect 2105 484 2109 553
rect 2112 532 2115 539
rect 2122 529 2126 560
rect 2150 553 2154 560
rect 2177 556 2181 560
rect 2192 563 2196 626
rect 2201 620 2229 623
rect 2208 614 2211 620
rect 2357 624 2382 627
rect 2392 627 2421 631
rect 2392 625 2398 627
rect 2357 622 2360 624
rect 2192 559 2209 563
rect 2217 562 2220 574
rect 2277 606 2287 609
rect 2232 569 2273 572
rect 2232 562 2235 569
rect 2238 562 2266 565
rect 2217 559 2235 562
rect 2221 556 2225 559
rect 2133 532 2136 549
rect 2143 549 2154 553
rect 2160 552 2225 556
rect 2245 556 2248 562
rect 2143 529 2147 549
rect 2150 532 2153 540
rect 2160 529 2164 552
rect 2177 505 2181 552
rect 2185 541 2213 544
rect 2192 535 2195 541
rect 2201 505 2204 515
rect 2216 532 2246 535
rect 2216 528 2219 532
rect 2238 531 2246 532
rect 2254 534 2257 546
rect 2270 534 2273 569
rect 2254 531 2273 534
rect 2277 528 2280 606
rect 2292 606 2302 609
rect 2310 609 2313 617
rect 2322 619 2360 622
rect 2392 621 2395 625
rect 2322 609 2325 619
rect 2363 618 2395 621
rect 2425 619 2434 623
rect 2363 615 2366 618
rect 2441 616 2445 638
rect 2449 627 2450 631
rect 2485 629 2488 638
rect 2529 629 2532 638
rect 2485 624 2497 629
rect 2529 624 2553 629
rect 2560 628 2564 638
rect 2595 628 2598 638
rect 2560 624 2587 628
rect 2595 625 2607 628
rect 2449 622 2457 624
rect 2454 619 2457 622
rect 2476 619 2477 623
rect 2485 616 2488 624
rect 2493 619 2501 624
rect 2520 619 2521 623
rect 2529 616 2532 624
rect 2560 623 2573 624
rect 2560 616 2564 623
rect 2595 620 2598 625
rect 2310 606 2325 609
rect 2310 603 2313 606
rect 2362 612 2368 615
rect 2301 593 2304 597
rect 2322 596 2327 599
rect 2340 599 2343 603
rect 2387 599 2390 603
rect 2433 606 2445 616
rect 2477 606 2488 616
rect 2521 606 2532 616
rect 2421 601 2425 606
rect 2457 601 2461 606
rect 2501 601 2505 606
rect 2552 601 2556 606
rect 2586 602 2589 610
rect 2332 596 2396 599
rect 2420 597 2564 601
rect 2579 599 2589 602
rect 2322 593 2325 596
rect 2295 590 2325 593
rect 2216 525 2280 528
rect 2216 505 2219 525
rect 2177 501 2193 505
rect 2201 502 2219 505
rect 2201 497 2204 502
rect 2299 498 2327 501
rect 2114 484 2118 489
rect 2135 484 2139 489
rect 2152 484 2156 489
rect 2300 492 2303 498
rect 2324 497 2327 498
rect 2324 494 2395 497
rect 2090 481 2157 484
rect 2192 479 2195 487
rect 2181 476 2195 479
rect 2281 468 2286 471
rect 2291 469 2301 472
rect 2309 472 2312 480
rect 2339 488 2342 494
rect 2358 488 2361 494
rect 2309 469 2330 472
rect 2309 466 2312 469
rect 2172 454 2175 461
rect 2172 451 2183 454
rect 2197 453 2201 461
rect 2237 454 2240 461
rect 2300 456 2303 460
rect 2231 451 2240 454
rect 2294 454 2318 456
rect 2294 453 2312 454
rect 2193 442 2211 445
rect 2167 434 2168 439
rect 2198 434 2201 442
rect 2156 420 2160 424
rect 2134 419 2137 420
rect 2033 416 2137 419
rect 2154 416 2160 420
rect 2167 416 2170 434
rect 1800 176 1805 187
rect 1832 181 1869 185
rect 1832 179 1836 181
rect 1659 170 1667 172
rect 1664 167 1667 170
rect 1686 167 1687 171
rect 1695 164 1698 172
rect 1703 167 1711 172
rect 1730 167 1731 171
rect 1739 164 1742 172
rect 1770 171 1805 176
rect 1815 175 1836 179
rect 1877 178 1880 187
rect 1909 183 1912 188
rect 1770 164 1774 171
rect 1643 154 1655 164
rect 1687 154 1698 164
rect 1731 154 1742 164
rect 1631 149 1635 154
rect 1667 149 1671 154
rect 1711 149 1715 154
rect 1762 149 1766 154
rect 1630 145 1774 149
rect 1634 119 1787 123
rect 1640 113 1644 119
rect 1678 113 1682 119
rect 1722 113 1726 119
rect 1767 113 1771 119
rect 1799 115 1804 171
rect 1815 127 1819 175
rect 1858 159 1861 165
rect 1900 159 1903 176
rect 1850 156 1903 159
rect 1843 142 1871 145
rect 1844 136 1847 142
rect 1868 141 1871 142
rect 1868 138 1939 141
rect 1815 125 1821 127
rect 1809 115 1827 116
rect 1690 88 1703 113
rect 1734 88 1747 113
rect 1799 112 1830 115
rect 1799 111 1827 112
rect 1835 113 1845 116
rect 1853 116 1856 124
rect 1883 132 1886 138
rect 1902 132 1905 138
rect 1853 113 1874 116
rect 1799 110 1811 111
rect 1853 110 1856 113
rect 1629 77 1636 81
rect 1640 69 1649 73
rect 1656 66 1660 88
rect 1664 77 1665 81
rect 1700 79 1703 88
rect 1744 79 1747 88
rect 1700 74 1712 79
rect 1744 74 1768 79
rect 1775 78 1779 88
rect 1817 78 1822 103
rect 1844 100 1847 104
rect 1838 98 1862 100
rect 1838 97 1856 98
rect 1861 97 1862 98
rect 1871 90 1874 113
rect 1912 132 1932 135
rect 1912 126 1915 132
rect 1929 126 1932 132
rect 1893 105 1896 108
rect 1893 102 1911 105
rect 2006 112 2009 188
rect 1921 95 1924 102
rect 1921 92 1938 95
rect 1843 89 1862 90
rect 1838 87 1862 89
rect 1871 87 1914 90
rect 1664 72 1672 74
rect 1669 69 1672 72
rect 1691 69 1692 73
rect 1700 66 1703 74
rect 1708 69 1716 74
rect 1735 69 1736 73
rect 1744 66 1747 74
rect 1775 73 1822 78
rect 1775 66 1779 73
rect 1648 56 1660 66
rect 1692 56 1703 66
rect 1736 56 1747 66
rect 1817 62 1822 73
rect 1844 81 1847 87
rect 1935 81 1938 92
rect 2006 85 2009 107
rect 2018 81 2022 186
rect 1900 76 1925 79
rect 1935 77 2022 81
rect 1900 74 1903 76
rect 1817 61 1827 62
rect 1817 58 1830 61
rect 1817 57 1827 58
rect 1835 58 1845 61
rect 1853 61 1856 69
rect 1865 71 1903 74
rect 1935 73 1938 77
rect 1865 61 1868 71
rect 1906 70 1938 73
rect 1906 67 1909 70
rect 1853 58 1868 61
rect 1636 51 1640 56
rect 1672 51 1676 56
rect 1716 51 1720 56
rect 1767 51 1771 56
rect 1853 55 1856 58
rect 1635 47 1779 51
rect 1905 64 1911 67
rect 1844 45 1847 49
rect 1865 48 1870 51
rect 1883 51 1886 55
rect 1930 51 1933 55
rect 1875 48 1939 51
rect 1865 45 1868 48
rect 1838 42 1868 45
rect 1983 20 2011 23
rect 1773 12 1926 16
rect 1949 15 1977 18
rect 1779 6 1783 12
rect 1817 6 1821 12
rect 1861 6 1865 12
rect 1906 6 1910 12
rect 1956 9 1959 15
rect 1990 14 1993 20
rect 1829 -19 1842 6
rect 1873 -19 1886 6
rect 1768 -30 1775 -26
rect 1779 -38 1788 -34
rect 1795 -41 1799 -19
rect 1803 -30 1804 -26
rect 1839 -28 1842 -19
rect 1883 -28 1886 -19
rect 1839 -33 1851 -28
rect 1883 -33 1907 -28
rect 1914 -29 1918 -19
rect 2018 1 2022 77
rect 2033 182 2038 416
rect 2093 377 2121 380
rect 2100 371 2103 377
rect 2136 359 2140 372
rect 2151 371 2156 372
rect 2169 371 2173 373
rect 2151 366 2173 371
rect 2177 371 2181 373
rect 2177 369 2183 371
rect 2197 369 2201 434
rect 2237 433 2240 451
rect 2317 453 2318 454
rect 2327 446 2330 469
rect 2368 488 2388 491
rect 2368 482 2371 488
rect 2385 482 2388 488
rect 2349 461 2352 464
rect 2349 458 2367 461
rect 2427 478 2580 482
rect 2433 472 2437 478
rect 2471 472 2475 478
rect 2515 472 2519 478
rect 2560 472 2564 478
rect 2586 473 2614 476
rect 2377 451 2380 458
rect 2377 448 2394 451
rect 2299 445 2318 446
rect 2294 443 2318 445
rect 2327 443 2370 446
rect 2300 437 2303 443
rect 2391 440 2394 448
rect 2483 447 2496 472
rect 2527 447 2540 472
rect 2593 467 2596 473
rect 2206 426 2234 429
rect 2213 420 2216 426
rect 2391 436 2429 440
rect 2356 432 2381 435
rect 2356 430 2359 432
rect 2177 366 2185 369
rect 2109 341 2112 351
rect 2121 341 2123 342
rect 2093 337 2101 341
rect 2109 338 2123 341
rect 2109 333 2112 338
rect 2130 335 2134 344
rect 2100 315 2103 323
rect 2093 312 2103 315
rect 2122 290 2126 295
rect 2137 290 2141 359
rect 2144 338 2147 345
rect 2154 335 2158 366
rect 2181 362 2185 366
rect 2197 365 2214 369
rect 2222 368 2225 380
rect 2237 375 2278 378
rect 2237 368 2240 375
rect 2243 368 2271 371
rect 2222 365 2240 368
rect 2226 362 2230 365
rect 2181 359 2230 362
rect 2165 338 2168 354
rect 2175 358 2230 359
rect 2250 362 2253 368
rect 2175 355 2188 358
rect 2175 335 2179 355
rect 2182 311 2186 355
rect 2190 347 2218 350
rect 2197 341 2200 347
rect 2206 311 2209 321
rect 2221 338 2251 341
rect 2221 323 2224 338
rect 2243 337 2251 338
rect 2259 340 2262 352
rect 2275 340 2278 375
rect 2259 337 2278 340
rect 2283 323 2286 417
rect 2291 414 2301 417
rect 2309 417 2312 425
rect 2321 427 2359 430
rect 2391 429 2394 436
rect 2321 417 2324 427
rect 2362 426 2394 429
rect 2433 428 2442 432
rect 2362 423 2365 426
rect 2449 425 2453 447
rect 2457 436 2458 440
rect 2493 438 2496 447
rect 2537 438 2540 447
rect 2493 433 2505 438
rect 2537 433 2561 438
rect 2568 437 2572 447
rect 2602 437 2605 447
rect 2568 433 2594 437
rect 2602 434 2614 437
rect 2457 431 2465 433
rect 2462 428 2465 431
rect 2484 428 2485 432
rect 2493 425 2496 433
rect 2501 428 2509 433
rect 2528 428 2529 432
rect 2537 425 2540 433
rect 2568 432 2581 433
rect 2568 425 2572 432
rect 2602 429 2605 434
rect 2309 414 2324 417
rect 2309 411 2312 414
rect 2361 420 2367 423
rect 2300 401 2303 405
rect 2321 404 2326 407
rect 2339 407 2342 411
rect 2386 407 2389 411
rect 2441 415 2453 425
rect 2485 415 2496 425
rect 2529 415 2540 425
rect 2429 410 2433 415
rect 2465 410 2469 415
rect 2509 410 2513 415
rect 2560 410 2564 415
rect 2593 411 2596 419
rect 2331 404 2395 407
rect 2428 406 2572 410
rect 2586 408 2596 411
rect 2321 401 2324 404
rect 2294 398 2324 401
rect 2221 320 2286 323
rect 2221 311 2224 320
rect 2182 307 2198 311
rect 2206 308 2224 311
rect 2206 303 2209 308
rect 2146 290 2150 295
rect 2167 290 2171 295
rect 2317 301 2345 304
rect 2318 295 2321 301
rect 2342 300 2345 301
rect 2342 297 2413 300
rect 2122 287 2181 290
rect 2197 285 2200 293
rect 2186 282 2200 285
rect 2294 271 2304 274
rect 2309 272 2319 275
rect 2327 275 2330 283
rect 2357 291 2360 297
rect 2376 291 2379 297
rect 2327 272 2348 275
rect 2327 269 2330 272
rect 2318 259 2321 263
rect 2312 257 2336 259
rect 2312 256 2330 257
rect 2335 256 2336 257
rect 2345 249 2348 272
rect 2386 291 2406 294
rect 2386 285 2389 291
rect 2403 285 2406 291
rect 2367 264 2370 267
rect 2367 261 2385 264
rect 2448 284 2601 288
rect 2454 278 2458 284
rect 2492 278 2496 284
rect 2536 278 2540 284
rect 2581 278 2585 284
rect 2609 279 2637 282
rect 2395 254 2398 261
rect 2395 251 2412 254
rect 2504 253 2517 278
rect 2548 253 2561 278
rect 2616 273 2619 279
rect 2317 248 2336 249
rect 2312 246 2336 248
rect 2345 246 2388 249
rect 2409 246 2412 251
rect 2318 240 2321 246
rect 2409 242 2450 246
rect 2374 235 2399 238
rect 2374 233 2377 235
rect 2174 216 2177 223
rect 2174 213 2185 216
rect 2199 215 2203 223
rect 2239 216 2242 223
rect 2233 213 2242 216
rect 2195 204 2213 207
rect 2200 195 2203 204
rect 2239 195 2242 213
rect 2285 217 2304 220
rect 2177 182 2182 186
rect 2033 179 2158 182
rect 2033 11 2038 179
rect 2155 178 2158 179
rect 2175 178 2182 182
rect 2112 140 2140 143
rect 2119 134 2122 140
rect 2157 125 2161 134
rect 2172 133 2177 134
rect 2172 128 2178 133
rect 2199 131 2203 195
rect 2208 188 2236 191
rect 2215 182 2218 188
rect 2152 121 2170 125
rect 2175 124 2179 128
rect 2199 127 2216 131
rect 2224 130 2227 142
rect 2239 137 2280 140
rect 2239 130 2242 137
rect 2245 130 2273 133
rect 2224 127 2242 130
rect 2228 124 2232 127
rect 2128 104 2131 114
rect 2140 104 2143 105
rect 2112 100 2120 104
rect 2128 101 2144 104
rect 2128 96 2131 101
rect 2140 100 2144 101
rect 2151 97 2155 106
rect 2119 78 2122 86
rect 2112 75 2122 78
rect 2143 52 2147 57
rect 2158 52 2162 121
rect 2175 120 2232 124
rect 2252 124 2255 130
rect 2165 100 2168 107
rect 2175 97 2179 120
rect 2184 73 2188 120
rect 2192 109 2220 112
rect 2199 103 2202 109
rect 2208 73 2211 83
rect 2223 100 2253 103
rect 2223 91 2226 100
rect 2245 99 2253 100
rect 2261 102 2264 114
rect 2277 102 2280 137
rect 2261 99 2280 102
rect 2285 91 2288 217
rect 2309 217 2319 220
rect 2327 220 2330 228
rect 2339 230 2377 233
rect 2409 232 2412 242
rect 2454 234 2463 238
rect 2339 220 2342 230
rect 2380 229 2412 232
rect 2470 231 2474 253
rect 2478 242 2479 246
rect 2514 244 2517 253
rect 2558 244 2561 253
rect 2514 239 2526 244
rect 2558 239 2582 244
rect 2589 243 2593 253
rect 2625 243 2628 253
rect 2589 239 2617 243
rect 2625 240 2637 243
rect 2478 237 2486 239
rect 2483 234 2486 237
rect 2505 234 2506 238
rect 2514 231 2517 239
rect 2522 234 2530 239
rect 2549 234 2550 238
rect 2558 231 2561 239
rect 2589 238 2602 239
rect 2589 231 2593 238
rect 2625 235 2628 240
rect 2380 226 2383 229
rect 2327 217 2342 220
rect 2327 214 2330 217
rect 2379 223 2385 226
rect 2462 221 2474 231
rect 2506 221 2517 231
rect 2550 221 2561 231
rect 2450 216 2454 221
rect 2486 216 2490 221
rect 2530 216 2534 221
rect 2581 216 2585 221
rect 2616 217 2619 225
rect 2318 204 2321 208
rect 2339 207 2344 210
rect 2357 210 2360 214
rect 2404 210 2407 214
rect 2449 212 2593 216
rect 2609 214 2619 217
rect 2349 207 2413 210
rect 2339 204 2342 207
rect 2312 201 2342 204
rect 2223 88 2288 91
rect 2223 73 2226 88
rect 2184 69 2200 73
rect 2208 70 2226 73
rect 2208 65 2211 70
rect 2167 52 2171 57
rect 2143 49 2185 52
rect 2199 47 2202 55
rect 2188 44 2202 47
rect 2078 27 2106 30
rect 2079 21 2082 27
rect 2103 26 2106 27
rect 2103 23 2174 26
rect 2028 1 2045 2
rect 2017 0 2059 1
rect 2017 -3 2065 0
rect 2070 -2 2080 1
rect 2088 1 2091 9
rect 2118 17 2121 23
rect 2137 17 2140 23
rect 2088 -2 2109 1
rect 2088 -5 2091 -2
rect 1914 -31 1927 -29
rect 1965 -31 1968 -21
rect 1999 -31 2002 -21
rect 2033 -31 2037 -11
rect 2079 -15 2082 -11
rect 2073 -17 2097 -15
rect 2073 -18 2091 -17
rect 2096 -18 2097 -17
rect 2106 -25 2109 -2
rect 2147 17 2167 20
rect 2147 11 2150 17
rect 2164 11 2167 17
rect 2210 16 2363 20
rect 2128 -10 2131 -7
rect 2128 -13 2146 -10
rect 2216 10 2220 16
rect 2254 10 2258 16
rect 2298 10 2302 16
rect 2343 10 2347 16
rect 2371 11 2399 14
rect 2156 -20 2159 -13
rect 2266 -15 2279 10
rect 2310 -15 2323 10
rect 2378 5 2381 11
rect 2156 -23 2173 -20
rect 2184 -23 2212 -22
rect 2078 -26 2097 -25
rect 2073 -28 2097 -26
rect 2106 -28 2149 -25
rect 2170 -26 2212 -23
rect 1803 -35 1811 -33
rect 1808 -38 1811 -35
rect 1830 -38 1831 -34
rect 1839 -41 1842 -33
rect 1847 -38 1855 -33
rect 1874 -38 1875 -34
rect 1883 -41 1886 -33
rect 1914 -34 1957 -31
rect 1914 -41 1918 -34
rect 1922 -35 1957 -34
rect 1965 -34 1991 -31
rect 1965 -39 1968 -34
rect 1982 -35 1991 -34
rect 1999 -34 2055 -31
rect 1999 -39 2002 -34
rect 2009 -35 2055 -34
rect 1787 -51 1799 -41
rect 1831 -51 1842 -41
rect 1875 -51 1886 -41
rect 1775 -56 1779 -51
rect 1811 -56 1815 -51
rect 1855 -56 1859 -51
rect 1906 -56 1910 -51
rect 1774 -60 1918 -56
rect 1956 -63 1959 -55
rect 1949 -66 1959 -63
rect 2051 -54 2055 -35
rect 2079 -34 2082 -28
rect 2170 -34 2173 -26
rect 2216 -34 2225 -30
rect 2135 -39 2160 -36
rect 2170 -38 2176 -34
rect 2232 -37 2236 -15
rect 2240 -26 2241 -22
rect 2276 -24 2279 -15
rect 2320 -24 2323 -15
rect 2276 -29 2288 -24
rect 2320 -29 2344 -24
rect 2351 -25 2355 -15
rect 2387 -25 2390 -15
rect 2351 -29 2379 -25
rect 2387 -28 2399 -25
rect 2240 -31 2248 -29
rect 2245 -34 2248 -31
rect 2267 -34 2268 -30
rect 2276 -37 2279 -29
rect 2284 -34 2292 -29
rect 2311 -34 2312 -30
rect 2320 -37 2323 -29
rect 2351 -30 2364 -29
rect 2351 -37 2355 -30
rect 2387 -33 2390 -28
rect 2135 -41 2138 -39
rect 2051 -57 2065 -54
rect 2070 -57 2080 -54
rect 2088 -54 2091 -46
rect 2100 -44 2138 -41
rect 2170 -42 2173 -38
rect 2100 -54 2103 -44
rect 2141 -45 2173 -42
rect 2141 -48 2144 -45
rect 2224 -47 2236 -37
rect 2268 -47 2279 -37
rect 2312 -47 2323 -37
rect 2088 -57 2103 -54
rect 1990 -66 1993 -58
rect 2088 -60 2091 -57
rect 1983 -69 1993 -66
rect 2140 -51 2146 -48
rect 2212 -52 2216 -47
rect 2248 -52 2252 -47
rect 2292 -52 2296 -47
rect 2343 -52 2347 -47
rect 2378 -51 2381 -43
rect 2211 -56 2355 -52
rect 2371 -54 2381 -51
rect 2079 -70 2082 -66
rect 2100 -67 2105 -64
rect 2118 -64 2121 -60
rect 2165 -64 2168 -60
rect 2110 -67 2174 -64
rect 2100 -70 2103 -67
rect 2073 -73 2103 -70
<< m2contact >>
rect 1965 865 1970 870
rect 1629 829 1634 834
rect 1659 837 1664 842
rect 1658 827 1663 832
rect 1686 829 1691 834
rect 1730 829 1735 834
rect 1813 755 1818 760
rect 1836 745 1841 750
rect 1813 738 1818 743
rect 1619 702 1624 707
rect 1649 710 1654 715
rect 1648 700 1653 705
rect 1676 702 1681 707
rect 1720 702 1725 707
rect 1941 711 1946 716
rect 1836 691 1841 696
rect 1981 856 1986 861
rect 1965 711 1970 717
rect 1957 666 1962 671
rect 1973 675 1978 680
rect 1964 654 1969 660
rect 1630 595 1635 600
rect 1660 603 1665 608
rect 1659 593 1664 598
rect 1687 595 1692 600
rect 1731 595 1736 600
rect 1998 845 2003 851
rect 1990 684 1995 689
rect 1981 636 1986 641
rect 1819 519 1824 524
rect 1834 510 1839 515
rect 1635 470 1640 475
rect 1665 478 1670 483
rect 1819 502 1824 507
rect 1664 468 1669 473
rect 1692 470 1697 475
rect 1736 470 1741 475
rect 1974 489 1979 494
rect 2018 837 2023 842
rect 2005 693 2010 698
rect 1997 627 2002 632
rect 1990 549 1995 554
rect 1834 456 1839 461
rect 1981 467 1986 472
rect 1632 376 1637 381
rect 1662 384 1667 389
rect 2168 865 2173 870
rect 2146 856 2151 861
rect 2121 845 2126 851
rect 2111 837 2116 842
rect 2018 617 2023 622
rect 2007 539 2012 544
rect 1998 434 2003 439
rect 1661 374 1666 379
rect 1689 376 1694 381
rect 1733 376 1738 381
rect 1989 353 1994 358
rect 1816 315 1821 320
rect 1831 307 1836 312
rect 1643 262 1648 267
rect 1673 270 1678 275
rect 1816 298 1821 303
rect 2017 424 2022 429
rect 2007 345 2012 350
rect 1672 260 1677 265
rect 1700 262 1705 267
rect 1744 262 1749 267
rect 1831 253 1836 258
rect 1996 261 2001 266
rect 1630 167 1635 172
rect 1660 175 1665 180
rect 2099 764 2104 769
rect 2118 764 2123 769
rect 2137 762 2142 767
rect 2155 764 2160 769
rect 2290 733 2295 738
rect 2320 741 2325 746
rect 2319 731 2324 736
rect 2347 733 2352 738
rect 2391 733 2396 738
rect 2274 657 2279 662
rect 2287 659 2292 664
rect 2152 636 2157 641
rect 2134 627 2139 632
rect 2123 617 2128 622
rect 2112 539 2117 544
rect 2131 549 2136 554
rect 2150 540 2155 545
rect 2287 605 2292 610
rect 2420 619 2425 624
rect 2450 627 2455 632
rect 2449 617 2454 622
rect 2477 619 2482 624
rect 2521 619 2526 624
rect 2276 466 2281 471
rect 2286 467 2291 472
rect 2168 434 2173 439
rect 2155 424 2160 429
rect 1659 165 1664 170
rect 1687 167 1692 172
rect 1731 167 1736 172
rect 1816 120 1821 125
rect 1830 111 1835 116
rect 1816 103 1821 108
rect 1635 69 1640 74
rect 1665 77 1670 82
rect 2018 186 2023 191
rect 2005 107 2010 112
rect 1664 67 1669 72
rect 1692 69 1697 74
rect 1736 69 1741 74
rect 1830 57 1835 62
rect 1774 -38 1779 -33
rect 1804 -30 1809 -25
rect 2144 345 2149 350
rect 2163 354 2168 359
rect 2286 413 2291 418
rect 2428 428 2433 433
rect 2458 436 2463 441
rect 2457 426 2462 431
rect 2485 428 2490 433
rect 2529 428 2534 433
rect 2289 269 2294 274
rect 2304 270 2309 275
rect 2177 186 2182 191
rect 2165 107 2170 112
rect 2304 216 2309 221
rect 2449 234 2454 239
rect 2479 242 2484 247
rect 2478 232 2483 237
rect 2506 234 2511 239
rect 2550 234 2555 239
rect 2033 6 2038 11
rect 2065 -4 2070 1
rect 2033 -11 2038 -6
rect 1803 -40 1808 -35
rect 1831 -38 1836 -33
rect 1875 -38 1880 -33
rect 2211 -34 2216 -29
rect 2241 -26 2246 -21
rect 2240 -36 2245 -31
rect 2268 -34 2273 -29
rect 2312 -34 2317 -29
rect 2065 -58 2070 -53
<< pm12contact >>
rect 1892 728 1897 733
rect 1901 727 1906 732
rect 1890 493 1895 498
rect 1899 492 1904 497
rect 1887 290 1892 295
rect 1896 289 1901 294
rect 2343 642 2348 647
rect 2352 641 2357 646
rect 1886 94 1891 99
rect 1895 93 1900 98
rect 2342 450 2347 455
rect 2351 449 2356 454
rect 2360 253 2365 258
rect 2369 252 2374 257
rect 2121 -21 2126 -16
rect 2130 -22 2135 -17
<< metal2 >>
rect 1659 887 1690 890
rect 1659 842 1663 887
rect 1686 834 1690 887
rect 1970 865 2168 870
rect 1986 856 2146 861
rect 2003 846 2121 851
rect 2023 837 2111 841
rect 1608 829 1629 833
rect 1620 805 1626 829
rect 1659 805 1663 827
rect 1730 805 1735 829
rect 1620 802 1739 805
rect 2320 791 2351 794
rect 2155 769 2160 770
rect 1649 760 1680 763
rect 1649 715 1653 760
rect 1676 707 1680 760
rect 1813 743 1818 755
rect 1837 739 1840 745
rect 1837 736 1874 739
rect 1871 733 1874 736
rect 1871 730 1892 733
rect 1901 717 1904 727
rect 1838 714 1904 717
rect 1598 702 1619 706
rect 1610 678 1616 702
rect 1649 678 1653 700
rect 1720 678 1725 702
rect 1838 696 1841 714
rect 1946 711 1965 716
rect 2099 698 2104 764
rect 2010 693 2104 698
rect 2118 689 2123 764
rect 1995 684 2123 689
rect 2137 680 2142 762
rect 1610 675 1729 678
rect 1978 675 2142 680
rect 2155 671 2160 764
rect 2320 746 2324 791
rect 2347 738 2351 791
rect 2269 733 2290 737
rect 2281 709 2287 733
rect 2320 709 2324 731
rect 2391 709 2396 733
rect 2281 706 2400 709
rect 1962 666 2160 671
rect 2450 677 2481 680
rect 2159 660 2274 662
rect 1660 653 1691 656
rect 1969 657 2274 660
rect 1969 655 2164 657
rect 1660 608 1664 653
rect 1687 600 1691 653
rect 2288 653 2291 659
rect 2288 650 2325 653
rect 2322 647 2325 650
rect 1986 636 2152 641
rect 2157 636 2158 641
rect 2322 644 2343 647
rect 2002 627 2134 632
rect 2139 627 2140 632
rect 2352 631 2355 641
rect 2289 628 2355 631
rect 2450 632 2454 677
rect 2023 618 2123 622
rect 2289 610 2292 628
rect 2477 624 2481 677
rect 2399 619 2420 623
rect 1609 595 1630 599
rect 1621 571 1627 595
rect 1660 571 1664 593
rect 1731 571 1736 595
rect 2411 595 2417 619
rect 2450 595 2454 617
rect 2521 595 2526 619
rect 2411 592 2530 595
rect 1621 568 1740 571
rect 1995 549 2131 554
rect 2012 539 2112 544
rect 1665 528 1696 531
rect 1665 483 1669 528
rect 1692 475 1696 528
rect 1819 507 1824 519
rect 1835 504 1838 510
rect 1835 501 1872 504
rect 1869 498 1872 501
rect 1869 495 1890 498
rect 2150 494 2155 540
rect 1899 482 1902 492
rect 1979 489 2155 494
rect 1836 479 1902 482
rect 2458 486 2489 489
rect 1614 470 1635 474
rect 1626 446 1632 470
rect 1665 446 1669 468
rect 1736 446 1741 470
rect 1836 461 1839 479
rect 1986 467 2276 471
rect 2287 461 2290 467
rect 2287 458 2324 461
rect 2321 455 2324 458
rect 1626 443 1745 446
rect 2321 452 2342 455
rect 2351 439 2354 449
rect 1662 434 1693 437
rect 2003 434 2168 439
rect 2288 436 2354 439
rect 2458 441 2462 486
rect 1662 389 1666 434
rect 1689 381 1693 434
rect 2022 424 2155 429
rect 2288 418 2291 436
rect 2485 433 2489 486
rect 2407 428 2428 432
rect 2419 404 2425 428
rect 2458 404 2462 426
rect 2529 404 2534 428
rect 2419 401 2538 404
rect 1611 376 1632 380
rect 1623 352 1629 376
rect 1662 352 1666 374
rect 1733 352 1738 376
rect 1988 358 2163 359
rect 1988 354 1989 358
rect 1994 354 2163 358
rect 1623 349 1742 352
rect 2012 345 2144 350
rect 1673 320 1704 323
rect 1673 275 1677 320
rect 1700 267 1704 320
rect 1816 303 1821 315
rect 1832 301 1835 307
rect 1832 298 1869 301
rect 1866 295 1869 298
rect 1866 292 1887 295
rect 2479 292 2510 295
rect 1896 279 1899 289
rect 1833 276 1899 279
rect 1622 262 1643 266
rect 1634 238 1640 262
rect 1673 238 1677 260
rect 1744 238 1749 262
rect 1833 258 1836 276
rect 2289 266 2294 269
rect 2001 261 2294 266
rect 2305 264 2308 270
rect 2305 261 2342 264
rect 2339 258 2342 261
rect 2339 255 2360 258
rect 2369 242 2372 252
rect 2479 247 2483 292
rect 2306 239 2372 242
rect 2506 239 2510 292
rect 1634 235 1753 238
rect 1660 225 1691 228
rect 1660 180 1664 225
rect 1687 172 1691 225
rect 2306 221 2309 239
rect 2428 234 2449 238
rect 2440 210 2446 234
rect 2479 210 2483 232
rect 2550 210 2555 234
rect 2440 207 2559 210
rect 2023 186 2177 191
rect 1609 167 1630 171
rect 1621 143 1627 167
rect 1660 143 1664 165
rect 1731 143 1736 167
rect 1621 140 1740 143
rect 1665 127 1696 130
rect 1665 82 1669 127
rect 1692 74 1696 127
rect 1816 108 1821 120
rect 1831 105 1834 111
rect 2010 107 2165 112
rect 1831 102 1868 105
rect 1865 99 1868 102
rect 1865 96 1886 99
rect 1895 83 1898 93
rect 1832 80 1898 83
rect 1614 69 1635 73
rect 1626 45 1632 69
rect 1665 45 1669 67
rect 1736 45 1741 69
rect 1832 62 1835 80
rect 1626 42 1745 45
rect 2241 24 2272 27
rect 1804 20 1835 23
rect 1804 -25 1808 20
rect 1831 -33 1835 20
rect 2033 -6 2038 6
rect 2066 -10 2069 -4
rect 2066 -13 2103 -10
rect 2100 -16 2103 -13
rect 2100 -19 2121 -16
rect 2241 -21 2245 24
rect 2130 -32 2133 -22
rect 2268 -29 2272 24
rect 1755 -38 1774 -34
rect 1765 -62 1771 -38
rect 1804 -62 1808 -40
rect 1875 -62 1880 -38
rect 2067 -35 2133 -32
rect 2190 -34 2211 -30
rect 2067 -53 2070 -35
rect 2202 -58 2208 -34
rect 2241 -58 2245 -36
rect 2312 -58 2317 -34
rect 2202 -61 2321 -58
rect 1765 -65 1884 -62
<< m123contact >>
rect 1844 776 1849 781
rect 1844 723 1849 728
rect 1862 727 1867 732
rect 1876 682 1881 687
rect 2295 690 2300 695
rect 2295 637 2300 642
rect 2313 641 2318 646
rect 2327 596 2332 601
rect 1842 541 1847 546
rect 1842 488 1847 493
rect 1860 492 1865 497
rect 2294 498 2299 503
rect 1874 447 1879 452
rect 2294 445 2299 450
rect 2312 449 2317 454
rect 2326 404 2331 409
rect 1839 338 1844 343
rect 2312 301 2317 306
rect 1839 285 1844 290
rect 1857 289 1862 294
rect 1871 244 1876 249
rect 2312 248 2317 253
rect 2330 252 2335 257
rect 2344 207 2349 212
rect 1838 142 1843 147
rect 1838 89 1843 94
rect 1856 93 1861 98
rect 1870 48 1875 53
rect 2073 27 2078 32
rect 2073 -26 2078 -21
rect 2091 -22 2096 -17
rect 2105 -67 2110 -62
<< metal3 >>
rect 1844 728 1847 776
rect 1867 727 1879 730
rect 1876 687 1879 727
rect 2295 642 2298 690
rect 2318 641 2330 644
rect 2327 601 2330 641
rect 1842 493 1845 541
rect 1865 492 1877 495
rect 1874 452 1877 492
rect 2294 450 2297 498
rect 2317 449 2329 452
rect 2326 409 2329 449
rect 1839 290 1842 338
rect 1862 289 1874 292
rect 1871 249 1874 289
rect 2312 253 2315 301
rect 2335 252 2347 255
rect 2344 212 2347 252
rect 1838 94 1841 142
rect 1861 93 1873 96
rect 1870 53 1873 93
rect 2073 -21 2076 27
rect 2096 -22 2108 -19
rect 2105 -62 2108 -22
<< labels >>
rlabel metal1 1862 676 1866 679 1 gnd
rlabel metal1 1912 682 1915 684 1 gnd
rlabel metal1 1860 732 1861 734 1 gnd
rlabel metal1 1856 776 1859 778 5 vdd
rlabel metal1 1857 722 1860 724 1 vdd
rlabel metal1 1833 746 1834 749 1 a3
rlabel metal1 1833 692 1834 695 1 b3
rlabel m2contact 1941 711 1945 715 7 p3
rlabel metal1 1919 835 1920 836 7 g3
rlabel metal1 1856 829 1857 830 3 b3
rlabel metal1 1855 836 1856 837 3 a3
rlabel metal1 1879 867 1879 867 5 vdd!
rlabel metal1 1879 803 1879 803 1 gnd!
rlabel metal1 1628 682 1631 683 1 gnd
rlabel metal1 1634 754 1636 755 5 vdd
rlabel metal2 1615 703 1615 703 1 clk_org
rlabel metal1 1618 711 1618 711 1 b3in
rlabel metal1 1769 710 1769 710 1 b3
rlabel metal1 1638 809 1641 810 1 gnd
rlabel metal1 1644 881 1646 882 5 vdd
rlabel metal2 1625 830 1625 830 1 clk_org
rlabel metal1 1626 839 1626 839 1 a3in
rlabel metal1 1780 835 1780 835 1 a3
rlabel metal1 1870 568 1870 568 1 gnd!
rlabel metal1 1870 632 1870 632 5 vdd!
rlabel metal1 1845 601 1846 602 3 a2
rlabel metal1 1847 594 1848 595 3 b2
rlabel metal1 1910 600 1911 601 7 g2
rlabel metal1 1939 476 1943 480 1 p2
rlabel metal1 1831 457 1832 460 1 b2
rlabel metal1 1831 511 1832 514 1 a2
rlabel metal1 1855 487 1858 489 1 vdd
rlabel metal1 1854 541 1857 543 5 vdd
rlabel metal1 1858 497 1859 499 1 gnd
rlabel metal1 1910 447 1913 449 1 gnd
rlabel metal1 1860 441 1864 444 1 gnd
rlabel metal1 1785 477 1785 477 1 b2
rlabel metal1 1633 480 1633 480 1 b2in
rlabel metal1 1779 602 1779 602 1 a2
rlabel metal1 1628 606 1628 606 1 a2in
rlabel metal2 1631 471 1631 471 1 clk_org
rlabel metal1 1650 522 1652 523 5 vdd
rlabel metal1 1644 450 1647 451 1 gnd
rlabel metal2 1626 596 1626 596 1 clk_org
rlabel metal1 1645 647 1647 648 5 vdd
rlabel metal1 1639 575 1642 576 1 gnd
rlabel metal1 1794 269 1794 269 1 b1
rlabel metal1 1641 272 1641 272 1 b1in
rlabel metal1 1781 382 1781 382 1 a1
rlabel metal1 1630 387 1630 387 1 a1in
rlabel metal2 1639 263 1639 263 1 clk_org
rlabel metal1 1658 314 1660 315 5 vdd
rlabel metal1 1652 242 1655 243 1 gnd
rlabel metal1 1641 356 1644 357 1 gnd
rlabel metal1 1647 428 1649 429 5 vdd
rlabel metal2 1628 377 1628 377 1 clk_org
rlabel metal1 1857 238 1861 241 1 gnd
rlabel metal1 1907 244 1910 246 1 gnd
rlabel metal1 1855 294 1856 296 1 gnd
rlabel metal1 1851 338 1854 340 5 vdd
rlabel metal1 1852 284 1855 286 1 vdd
rlabel metal1 1828 254 1829 257 1 b1
rlabel metal1 1828 308 1829 311 1 a1
rlabel space 1936 273 1940 277 1 p1
rlabel metal1 1878 349 1878 349 1 gnd!
rlabel metal1 1878 413 1878 413 5 vdd!
rlabel metal1 1854 382 1855 383 3 a1
rlabel metal1 1855 375 1856 376 3 b1
rlabel metal1 1918 381 1919 382 7 g1
rlabel metal2 1626 168 1626 168 1 clk_org
rlabel metal1 1645 219 1647 220 5 vdd
rlabel metal1 1639 147 1642 148 1 gnd
rlabel metal2 1631 70 1631 70 1 clk_org
rlabel metal1 1650 121 1652 122 5 vdd
rlabel metal1 1644 49 1647 50 1 gnd
rlabel metal1 1629 177 1629 177 1 a0in
rlabel metal1 1778 174 1778 174 1 a0
rlabel metal1 1632 79 1632 79 1 b0in
rlabel metal1 1785 76 1785 76 1 b0
rlabel metal1 1827 58 1828 61 1 b0
rlabel metal1 1827 112 1828 115 1 a0
rlabel metal1 1935 77 1939 81 7 p0
rlabel metal1 1851 88 1854 90 1 vdd
rlabel metal1 1850 142 1853 144 5 vdd
rlabel metal1 1854 98 1855 100 1 gnd
rlabel metal1 1906 48 1909 50 1 gnd
rlabel metal1 1856 42 1860 45 1 gnd
rlabel metal1 1876 221 1876 221 5 vdd!
rlabel metal1 1876 157 1876 157 1 gnd!
rlabel metal1 1851 190 1852 191 3 a0
rlabel metal1 1853 183 1854 184 3 b0
rlabel metal1 1916 189 1917 190 7 g0
rlabel metal2 1770 -37 1770 -37 1 clk_org
rlabel metal1 1789 14 1791 15 5 vdd
rlabel metal1 1783 -58 1786 -57 1 gnd
rlabel metal1 1769 -28 1769 -28 1 cinin
rlabel metal1 2173 833 2174 834 1 p3
rlabel metal1 2150 833 2151 834 1 p2
rlabel metal1 2123 833 2124 834 1 p1
rlabel metal1 2156 756 2157 757 1 g3
rlabel metal1 2121 755 2122 756 1 g1
rlabel metal1 2100 755 2101 756 1 g0
rlabel metal1 2189 699 2191 700 1 gnd
rlabel metal1 2197 764 2199 765 1 vdd
rlabel metal1 2111 833 2112 835 1 p0
rlabel metal1 2255 785 2262 786 1 vdd
rlabel metal1 2218 843 2225 844 1 vdd
rlabel metal1 2205 781 2211 785 1 clk
rlabel metal1 2220 724 2223 757 1 c3
rlabel metal1 2182 831 2193 835 1 c3bar
rlabel metal1 2075 754 2078 758 3 clk
rlabel metal1 2085 751 2089 760 1 gnd
rlabel metal1 2063 755 2075 758 1 clk
rlabel metal1 2047 754 2055 758 1 clk_org
rlabel metal1 2047 730 2049 731 1 gnd
rlabel metal1 2055 795 2057 796 1 vdd
rlabel metal1 2138 755 2139 756 1 g2
rlabel metal1 2197 860 2200 872 3 clk
rlabel metal1 2196 880 2200 888 3 clk_org
rlabel metal1 2172 886 2173 888 3 gnd
rlabel metal1 2237 878 2238 880 3 vdd
rlabel metal1 2233 644 2234 646 3 vdd
rlabel metal1 2168 652 2169 654 3 gnd
rlabel metal1 2192 646 2196 654 3 clk_org
rlabel metal1 2193 626 2196 638 3 clk
rlabel metal1 2068 572 2070 573 1 vdd
rlabel metal1 2060 507 2062 508 1 gnd
rlabel metal1 2060 531 2068 535 1 clk_org
rlabel metal1 2076 532 2088 535 1 clk
rlabel metal1 2216 502 2219 535 1 c2
rlabel metal1 2177 501 2181 565 1 c2bar
rlabel metal1 2098 529 2102 538 1 gnd
rlabel metal1 2088 532 2091 536 3 clk
rlabel metal1 2124 611 2125 613 1 p0
rlabel metal1 2113 533 2114 534 1 g0
rlabel metal1 2134 533 2135 534 1 g1
rlabel metal1 2151 533 2152 534 1 g2
rlabel metal1 2136 611 2137 612 1 p1
rlabel metal1 2163 611 2164 612 1 p2
rlabel metal1 2201 559 2207 563 1 clk
rlabel metal1 2214 621 2221 622 1 vdd
rlabel metal1 2251 563 2258 564 1 vdd
rlabel metal1 2193 542 2195 543 1 vdd
rlabel metal1 2185 477 2187 478 1 gnd
rlabel metal1 2284 606 2285 609 1 c2
rlabel metal1 2313 590 2317 593 1 gnd
rlabel metal1 2363 596 2366 598 1 gnd
rlabel metal1 2311 646 2312 648 1 gnd
rlabel metal1 2307 690 2310 692 5 vdd
rlabel metal1 2308 636 2311 638 1 vdd
rlabel metal1 2284 660 2285 663 1 p3
rlabel metal1 2101 378 2103 379 1 vdd
rlabel metal1 2093 313 2095 314 1 gnd
rlabel metal1 2093 337 2101 341 1 clk_org
rlabel metal1 2109 338 2121 341 1 clk
rlabel metal1 2198 433 2201 445 3 clk
rlabel metal1 2197 453 2201 461 3 clk_org
rlabel metal1 2173 459 2174 461 3 gnd
rlabel metal1 2238 451 2239 453 3 vdd
rlabel metal1 2221 308 2224 341 1 c1
rlabel metal1 2181 355 2188 362 1 c1bar
rlabel metal1 2168 417 2169 418 1 p1
rlabel metal1 2166 339 2167 340 1 g1
rlabel metal1 2145 339 2146 340 1 g0
rlabel metal1 2156 417 2157 419 1 p0
rlabel space 2120 338 2123 342 3 clk
rlabel metal1 2130 335 2134 344 1 gnd
rlabel metal1 2206 365 2212 369 1 clk
rlabel metal1 2219 427 2226 428 1 vdd
rlabel metal1 2256 369 2263 370 1 vdd
rlabel metal1 2198 348 2200 349 1 vdd
rlabel metal1 2190 283 2192 284 1 gnd
rlabel metal1 2128 101 2140 104 1 clk
rlabel metal1 2112 100 2120 104 1 clk_org
rlabel metal1 2112 76 2114 77 1 gnd
rlabel metal1 2120 141 2122 142 1 vdd
rlabel metal1 2240 213 2241 215 3 vdd
rlabel metal1 2175 221 2176 223 3 gnd
rlabel metal1 2199 215 2203 223 3 clk_org
rlabel metal1 2200 195 2203 207 3 clk
rlabel metal1 2223 70 2226 103 1 c0
rlabel metal1 2175 120 2232 124 1 c0bar
rlabel metal1 2166 101 2167 102 1 g0
rlabel metal1 2177 179 2178 181 1 p0
rlabel metal1 2141 100 2144 104 3 clk
rlabel metal1 2151 97 2155 106 1 gnd
rlabel metal1 2208 127 2214 131 1 clk
rlabel metal1 2221 189 2228 190 1 vdd
rlabel metal1 2258 131 2265 132 1 vdd
rlabel metal1 2200 110 2202 111 1 vdd
rlabel metal1 2192 45 2194 46 1 gnd
rlabel metal1 2330 201 2334 204 1 gnd
rlabel metal1 2380 207 2383 209 1 gnd
rlabel metal1 2324 301 2327 303 5 vdd
rlabel metal1 2325 247 2328 249 1 vdd
rlabel metal1 2301 271 2302 274 1 p1
rlabel metal1 2328 257 2329 259 1 gnd
rlabel metal1 2301 217 2302 220 1 c0
rlabel metal1 2458 214 2461 215 1 gnd
rlabel metal1 2464 286 2466 287 5 vdd
rlabel metal2 2445 235 2445 235 1 clk_org
rlabel metal1 2448 243 2448 243 1 s1in
rlabel metal1 2599 240 2599 240 1 s1
rlabel metal1 2613 240 2613 240 1 s1
rlabel metal1 2609 215 2611 216 1 gnd
rlabel metal1 2617 280 2619 281 1 vdd
rlabel metal1 2429 599 2432 600 1 gnd
rlabel metal1 2435 671 2437 672 5 vdd
rlabel metal2 2416 620 2416 620 1 clk_org
rlabel metal1 2417 628 2417 628 1 s3in
rlabel metal1 2570 625 2570 625 1 s3
rlabel metal1 2586 625 2586 625 1 s3
rlabel metal1 2579 600 2581 601 1 gnd
rlabel metal1 2587 665 2589 666 1 vdd
rlabel metal1 2440 739 2440 739 7 cout
rlabel metal1 2287 743 2287 743 1 c3
rlabel metal2 2286 734 2286 734 1 clk_org
rlabel metal1 2305 785 2307 786 5 vdd
rlabel metal1 2299 713 2302 714 1 gnd
rlabel metal1 2457 778 2459 779 1 vdd
rlabel metal1 2449 713 2451 714 1 gnd
rlabel metal1 2452 738 2452 738 1 cout
rlabel metal1 2589 434 2589 434 1 s2
rlabel metal1 2586 409 2588 410 1 gnd
rlabel metal1 2594 474 2596 475 1 vdd
rlabel metal1 2577 435 2577 435 1 s2
rlabel metal1 2425 438 2425 438 1 s2in
rlabel metal2 2424 429 2424 429 1 clk_org
rlabel metal1 2443 480 2445 481 5 vdd
rlabel metal1 2437 408 2440 409 1 gnd
rlabel metal1 2283 414 2284 417 1 c1
rlabel metal1 2283 468 2284 471 1 p2
rlabel metal1 2307 444 2310 446 1 vdd
rlabel metal1 2306 498 2309 500 5 vdd
rlabel metal1 2310 454 2311 456 1 gnd
rlabel metal1 2362 404 2365 406 1 gnd
rlabel metal1 2312 398 2316 401 1 gnd
rlabel metal1 2174 -36 2174 -36 1 s0in
rlabel metal1 2062 -3 2063 0 1 p0
rlabel metal1 2086 -27 2089 -25 1 vdd
rlabel metal1 2085 27 2088 29 5 vdd
rlabel metal1 2089 -17 2090 -15 1 gnd
rlabel metal1 2141 -67 2144 -65 1 gnd
rlabel metal1 2091 -73 2095 -70 1 gnd
rlabel metal1 2062 -55 2062 -55 1 cin2
rlabel metal1 1952 -33 1952 -33 1 cin
rlabel metal1 1957 16 1959 17 1 vdd
rlabel metal1 1949 -65 1951 -64 1 gnd
rlabel metal1 1974 -32 1974 -32 1 cin1
rlabel metal1 2009 -33 2009 -33 1 cin2
rlabel metal1 1985 -34 1985 -34 1 cin1
rlabel metal1 1991 21 1993 22 1 vdd
rlabel metal1 1983 -68 1985 -67 1 gnd
rlabel metal1 1924 -34 1924 -34 1 cin
rlabel metal1 2157 179 2157 179 1 cin2
rlabel metal1 2135 417 2135 417 1 cin2
rlabel metal1 2102 612 2102 612 1 cin2
rlabel metal1 2090 834 2090 834 1 cin2
rlabel metal1 2379 12 2381 13 1 vdd
rlabel metal1 2371 -53 2373 -52 1 gnd
rlabel metal2 2207 -33 2207 -33 1 clk_org
rlabel metal1 2226 18 2228 19 5 vdd
rlabel metal1 2220 -54 2223 -53 1 gnd
rlabel metal1 2287 -29 2287 -29 1 x
rlabel metal1 2330 -26 2330 -26 1 y
rlabel metal1 2365 -27 2365 -27 1 s0
<< end >>
