magic
tech scmos
timestamp 1732021615
<< nwell >>
rect 806 1091 830 1115
rect 845 1105 879 1111
rect 845 1075 907 1105
rect 946 1091 970 1115
rect 985 1105 1019 1111
rect 985 1075 1047 1105
rect 1081 1091 1105 1115
rect 1120 1105 1154 1111
rect 1120 1075 1182 1105
rect 1219 1090 1243 1114
rect 1258 1104 1292 1110
rect 873 1069 907 1075
rect 1013 1069 1047 1075
rect 1148 1069 1182 1075
rect 1258 1074 1320 1104
rect 1286 1068 1320 1074
rect 806 1036 830 1060
rect 946 1036 970 1060
rect 1081 1036 1105 1060
rect 1219 1035 1243 1059
rect 483 983 515 1020
rect 521 983 547 1020
rect 565 983 591 1020
rect 610 983 636 1020
rect 731 964 768 990
rect 774 964 802 990
rect 996 943 1024 977
rect 1168 964 1192 988
rect 1207 978 1241 984
rect 1207 948 1269 978
rect 1235 942 1269 948
rect 487 885 519 922
rect 525 885 551 922
rect 569 885 595 922
rect 614 885 640 922
rect 731 890 768 916
rect 774 890 802 916
rect 1168 909 1192 933
rect 1026 853 1054 907
rect 1368 889 1400 926
rect 1406 889 1432 926
rect 1450 889 1476 926
rect 1495 889 1521 926
rect 1574 891 1602 925
rect 492 787 524 824
rect 530 787 556 824
rect 574 787 600 824
rect 619 787 645 824
rect 731 821 768 847
rect 774 821 802 847
rect 1010 794 1038 828
rect 1063 825 1091 849
rect 1366 789 1398 826
rect 1404 789 1430 826
rect 1448 789 1474 826
rect 1493 789 1519 826
rect 1578 788 1606 822
rect 731 747 768 773
rect 774 747 802 773
rect 499 687 531 724
rect 537 687 563 724
rect 581 687 607 724
rect 626 687 652 724
rect 992 705 1020 739
rect 1166 731 1190 755
rect 1205 745 1239 751
rect 1205 715 1267 745
rect 1233 709 1267 715
rect 1166 676 1190 700
rect 1365 682 1397 719
rect 1403 682 1429 719
rect 1447 682 1473 719
rect 1492 682 1518 719
rect 1580 689 1608 723
rect 1022 615 1050 669
rect 510 573 542 610
rect 548 573 574 610
rect 592 573 618 610
rect 637 573 663 610
rect 1006 556 1034 590
rect 1059 587 1087 611
rect 1169 607 1193 631
rect 1208 621 1242 627
rect 1208 591 1270 621
rect 1236 585 1270 591
rect 1365 578 1397 615
rect 1403 578 1429 615
rect 1447 578 1473 615
rect 1492 578 1518 615
rect 1576 587 1604 621
rect 1169 552 1193 576
rect 502 464 534 501
rect 540 464 566 501
rect 584 464 610 501
rect 629 464 655 501
rect 997 478 1025 512
rect 1163 459 1187 483
rect 1202 473 1236 479
rect 1202 443 1264 473
rect 1365 463 1397 500
rect 1403 463 1429 500
rect 1447 463 1473 500
rect 1492 463 1518 500
rect 1573 468 1601 502
rect 1027 388 1055 442
rect 1230 437 1264 443
rect 1163 404 1187 428
rect 507 339 539 376
rect 545 339 571 376
rect 589 339 615 376
rect 634 339 660 376
rect 1011 329 1039 363
rect 1064 360 1092 384
rect 523 228 555 265
rect 561 228 587 265
rect 605 228 631 265
rect 650 228 676 265
rect 999 255 1027 289
rect 1029 165 1057 219
rect 513 110 545 147
rect 551 110 577 147
rect 595 110 621 147
rect 640 110 666 147
rect 1013 106 1041 140
rect 1066 137 1094 161
<< ntransistor >>
rect 817 1077 819 1083
rect 957 1077 959 1083
rect 1092 1077 1094 1083
rect 856 1028 858 1040
rect 866 1028 868 1040
rect 884 1028 886 1040
rect 894 1028 896 1040
rect 1230 1076 1232 1082
rect 996 1028 998 1040
rect 1006 1028 1008 1040
rect 1024 1028 1026 1040
rect 1034 1028 1036 1040
rect 1131 1028 1133 1040
rect 1141 1028 1143 1040
rect 1159 1028 1161 1040
rect 1169 1028 1171 1040
rect 817 1022 819 1028
rect 957 1022 959 1028
rect 1092 1022 1094 1028
rect 1269 1027 1271 1039
rect 1279 1027 1281 1039
rect 1297 1027 1299 1039
rect 1307 1027 1309 1039
rect 1230 1021 1232 1027
rect 490 957 492 967
rect 526 957 528 967
rect 534 957 536 967
rect 570 957 572 967
rect 578 957 580 967
rect 621 957 623 967
rect 744 936 746 949
rect 754 936 756 949
rect 786 947 788 954
rect 1179 950 1181 956
rect 1008 923 1010 933
rect 1218 901 1220 913
rect 1228 901 1230 913
rect 1246 901 1248 913
rect 1256 901 1258 913
rect 494 859 496 869
rect 530 859 532 869
rect 538 859 540 869
rect 574 859 576 869
rect 582 859 584 869
rect 625 859 627 869
rect 744 862 746 875
rect 754 862 756 875
rect 786 873 788 880
rect 917 853 919 894
rect 924 853 926 894
rect 950 854 952 894
rect 977 854 979 894
rect 1000 854 1002 894
rect 1179 895 1181 901
rect 1375 863 1377 873
rect 1411 863 1413 873
rect 1419 863 1421 873
rect 1455 863 1457 873
rect 1463 863 1465 873
rect 1506 863 1508 873
rect 1586 871 1588 881
rect 744 793 746 806
rect 754 793 756 806
rect 786 804 788 811
rect 903 776 905 816
rect 927 776 929 816
rect 948 776 950 816
rect 965 776 967 816
rect 983 777 985 817
rect 1022 774 1024 784
rect 499 761 501 771
rect 535 761 537 771
rect 543 761 545 771
rect 579 761 581 771
rect 587 761 589 771
rect 630 761 632 771
rect 1373 763 1375 773
rect 1409 763 1411 773
rect 1417 763 1419 773
rect 1453 763 1455 773
rect 1461 763 1463 773
rect 1504 763 1506 773
rect 1590 768 1592 778
rect 744 719 746 732
rect 754 719 756 732
rect 786 730 788 737
rect 1177 717 1179 723
rect 1004 685 1006 695
rect 506 661 508 671
rect 542 661 544 671
rect 550 661 552 671
rect 586 661 588 671
rect 594 661 596 671
rect 637 661 639 671
rect 1216 668 1218 680
rect 1226 668 1228 680
rect 1244 668 1246 680
rect 1254 668 1256 680
rect 930 615 932 656
rect 937 615 939 656
rect 963 616 965 656
rect 990 616 992 656
rect 1177 662 1179 668
rect 1592 669 1594 679
rect 1372 656 1374 666
rect 1408 656 1410 666
rect 1416 656 1418 666
rect 1452 656 1454 666
rect 1460 656 1462 666
rect 1503 656 1505 666
rect 517 547 519 557
rect 553 547 555 557
rect 561 547 563 557
rect 597 547 599 557
rect 605 547 607 557
rect 648 547 650 557
rect 916 538 918 578
rect 940 538 942 578
rect 961 538 963 578
rect 978 538 980 578
rect 1180 593 1182 599
rect 1018 536 1020 546
rect 1588 567 1590 577
rect 1219 544 1221 556
rect 1229 544 1231 556
rect 1247 544 1249 556
rect 1257 544 1259 556
rect 1372 552 1374 562
rect 1408 552 1410 562
rect 1416 552 1418 562
rect 1452 552 1454 562
rect 1460 552 1462 562
rect 1503 552 1505 562
rect 1180 538 1182 544
rect 1009 458 1011 468
rect 509 438 511 448
rect 545 438 547 448
rect 553 438 555 448
rect 589 438 591 448
rect 597 438 599 448
rect 640 438 642 448
rect 1174 445 1176 451
rect 962 388 964 429
rect 969 388 971 429
rect 995 389 997 429
rect 1585 448 1587 458
rect 1372 437 1374 447
rect 1408 437 1410 447
rect 1416 437 1418 447
rect 1452 437 1454 447
rect 1460 437 1462 447
rect 1503 437 1505 447
rect 1213 396 1215 408
rect 1223 396 1225 408
rect 1241 396 1243 408
rect 1251 396 1253 408
rect 1174 390 1176 396
rect 514 313 516 323
rect 550 313 552 323
rect 558 313 560 323
rect 594 313 596 323
rect 602 313 604 323
rect 645 313 647 323
rect 948 311 950 351
rect 972 311 974 351
rect 993 311 995 351
rect 1023 309 1025 319
rect 1011 235 1013 245
rect 530 202 532 212
rect 566 202 568 212
rect 574 202 576 212
rect 610 202 612 212
rect 618 202 620 212
rect 661 202 663 212
rect 983 165 985 206
rect 990 165 992 206
rect 520 84 522 94
rect 556 84 558 94
rect 564 84 566 94
rect 600 84 602 94
rect 608 84 610 94
rect 651 84 653 94
rect 969 88 971 128
rect 993 88 995 128
rect 1025 86 1027 96
<< ptransistor >>
rect 817 1097 819 1109
rect 856 1081 858 1105
rect 866 1081 868 1105
rect 884 1075 886 1099
rect 894 1075 896 1099
rect 957 1097 959 1109
rect 996 1081 998 1105
rect 1006 1081 1008 1105
rect 817 1042 819 1054
rect 1024 1075 1026 1099
rect 1034 1075 1036 1099
rect 1092 1097 1094 1109
rect 1131 1081 1133 1105
rect 1141 1081 1143 1105
rect 957 1042 959 1054
rect 1159 1075 1161 1099
rect 1169 1075 1171 1099
rect 1230 1096 1232 1108
rect 1269 1080 1271 1104
rect 1279 1080 1281 1104
rect 1092 1042 1094 1054
rect 1297 1074 1299 1098
rect 1307 1074 1309 1098
rect 1230 1041 1232 1053
rect 494 989 496 1014
rect 502 989 504 1014
rect 532 989 534 1014
rect 576 989 578 1014
rect 621 989 623 1014
rect 744 972 746 984
rect 754 972 756 984
rect 786 972 788 984
rect 1008 951 1010 971
rect 1179 970 1181 982
rect 1218 954 1220 978
rect 1228 954 1230 978
rect 1246 948 1248 972
rect 1256 948 1258 972
rect 498 891 500 916
rect 506 891 508 916
rect 536 891 538 916
rect 580 891 582 916
rect 625 891 627 916
rect 1179 915 1181 927
rect 744 898 746 910
rect 754 898 756 910
rect 786 898 788 910
rect 1038 861 1040 901
rect 1379 895 1381 920
rect 1387 895 1389 920
rect 1417 895 1419 920
rect 1461 895 1463 920
rect 1506 895 1508 920
rect 1586 899 1588 919
rect 744 829 746 841
rect 754 829 756 841
rect 786 829 788 841
rect 1075 833 1077 843
rect 503 793 505 818
rect 511 793 513 818
rect 541 793 543 818
rect 585 793 587 818
rect 630 793 632 818
rect 1022 802 1024 822
rect 1377 795 1379 820
rect 1385 795 1387 820
rect 1415 795 1417 820
rect 1459 795 1461 820
rect 1504 795 1506 820
rect 1590 796 1592 816
rect 744 755 746 767
rect 754 755 756 767
rect 786 755 788 767
rect 1177 737 1179 749
rect 510 693 512 718
rect 518 693 520 718
rect 548 693 550 718
rect 592 693 594 718
rect 637 693 639 718
rect 1004 713 1006 733
rect 1216 721 1218 745
rect 1226 721 1228 745
rect 1244 715 1246 739
rect 1254 715 1256 739
rect 1177 682 1179 694
rect 1376 688 1378 713
rect 1384 688 1386 713
rect 1414 688 1416 713
rect 1458 688 1460 713
rect 1503 688 1505 713
rect 1592 697 1594 717
rect 1034 623 1036 663
rect 1180 613 1182 625
rect 521 579 523 604
rect 529 579 531 604
rect 559 579 561 604
rect 603 579 605 604
rect 648 579 650 604
rect 1071 595 1073 605
rect 1018 564 1020 584
rect 1219 597 1221 621
rect 1229 597 1231 621
rect 1247 591 1249 615
rect 1257 591 1259 615
rect 1180 558 1182 570
rect 1376 584 1378 609
rect 1384 584 1386 609
rect 1414 584 1416 609
rect 1458 584 1460 609
rect 1503 584 1505 609
rect 1588 595 1590 615
rect 513 470 515 495
rect 521 470 523 495
rect 551 470 553 495
rect 595 470 597 495
rect 640 470 642 495
rect 1009 486 1011 506
rect 1174 465 1176 477
rect 1213 449 1215 473
rect 1223 449 1225 473
rect 1376 469 1378 494
rect 1384 469 1386 494
rect 1414 469 1416 494
rect 1458 469 1460 494
rect 1503 469 1505 494
rect 1585 476 1587 496
rect 1039 396 1041 436
rect 1241 443 1243 467
rect 1251 443 1253 467
rect 1174 410 1176 422
rect 518 345 520 370
rect 526 345 528 370
rect 556 345 558 370
rect 600 345 602 370
rect 645 345 647 370
rect 1076 368 1078 378
rect 1023 337 1025 357
rect 1011 263 1013 283
rect 534 234 536 259
rect 542 234 544 259
rect 572 234 574 259
rect 616 234 618 259
rect 661 234 663 259
rect 1041 173 1043 213
rect 1078 145 1080 155
rect 524 116 526 141
rect 532 116 534 141
rect 562 116 564 141
rect 606 116 608 141
rect 651 116 653 141
rect 1025 114 1027 134
<< ndiffusion >>
rect 816 1077 817 1083
rect 819 1077 820 1083
rect 956 1077 957 1083
rect 959 1077 960 1083
rect 1091 1077 1092 1083
rect 1094 1077 1095 1083
rect 855 1028 856 1040
rect 858 1028 866 1040
rect 868 1028 869 1040
rect 883 1028 884 1040
rect 886 1028 894 1040
rect 896 1028 897 1040
rect 1229 1076 1230 1082
rect 1232 1076 1233 1082
rect 995 1028 996 1040
rect 998 1028 1006 1040
rect 1008 1028 1009 1040
rect 1023 1028 1024 1040
rect 1026 1028 1034 1040
rect 1036 1028 1037 1040
rect 1130 1028 1131 1040
rect 1133 1028 1141 1040
rect 1143 1028 1144 1040
rect 1158 1028 1159 1040
rect 1161 1028 1169 1040
rect 1171 1028 1172 1040
rect 816 1022 817 1028
rect 819 1022 820 1028
rect 956 1022 957 1028
rect 959 1022 960 1028
rect 1091 1022 1092 1028
rect 1094 1022 1095 1028
rect 1268 1027 1269 1039
rect 1271 1027 1279 1039
rect 1281 1027 1282 1039
rect 1296 1027 1297 1039
rect 1299 1027 1307 1039
rect 1309 1027 1310 1039
rect 1229 1021 1230 1027
rect 1232 1021 1233 1027
rect 489 957 490 967
rect 492 957 493 967
rect 525 957 526 967
rect 528 957 529 967
rect 533 957 534 967
rect 536 957 537 967
rect 569 957 570 967
rect 572 957 573 967
rect 577 957 578 967
rect 580 957 581 967
rect 620 957 621 967
rect 623 957 624 967
rect 743 936 744 949
rect 746 936 754 949
rect 756 936 757 949
rect 785 947 786 954
rect 788 947 789 954
rect 1178 950 1179 956
rect 1181 950 1182 956
rect 1007 923 1008 933
rect 1010 923 1011 933
rect 1217 901 1218 913
rect 1220 901 1228 913
rect 1230 901 1231 913
rect 1245 901 1246 913
rect 1248 901 1256 913
rect 1258 901 1259 913
rect 493 859 494 869
rect 496 859 497 869
rect 529 859 530 869
rect 532 859 533 869
rect 537 859 538 869
rect 540 859 541 869
rect 573 859 574 869
rect 576 859 577 869
rect 581 859 582 869
rect 584 859 585 869
rect 624 859 625 869
rect 627 859 628 869
rect 743 862 744 875
rect 746 862 754 875
rect 756 862 757 875
rect 785 873 786 880
rect 788 873 789 880
rect 916 853 917 894
rect 919 853 924 894
rect 926 853 927 894
rect 949 854 950 894
rect 952 854 953 894
rect 976 854 977 894
rect 979 854 980 894
rect 999 854 1000 894
rect 1002 854 1003 894
rect 1178 895 1179 901
rect 1181 895 1182 901
rect 1374 863 1375 873
rect 1377 863 1378 873
rect 1410 863 1411 873
rect 1413 863 1414 873
rect 1418 863 1419 873
rect 1421 863 1422 873
rect 1454 863 1455 873
rect 1457 863 1458 873
rect 1462 863 1463 873
rect 1465 863 1466 873
rect 1505 863 1506 873
rect 1508 863 1509 873
rect 1585 871 1586 881
rect 1588 871 1589 881
rect 743 793 744 806
rect 746 793 754 806
rect 756 793 757 806
rect 785 804 786 811
rect 788 804 789 811
rect 902 776 903 816
rect 905 776 906 816
rect 926 776 927 816
rect 929 776 930 816
rect 947 776 948 816
rect 950 776 951 816
rect 964 776 965 816
rect 967 776 968 816
rect 982 777 983 817
rect 985 777 986 817
rect 1021 774 1022 784
rect 1024 774 1025 784
rect 498 761 499 771
rect 501 761 502 771
rect 534 761 535 771
rect 537 761 538 771
rect 542 761 543 771
rect 545 761 546 771
rect 578 761 579 771
rect 581 761 582 771
rect 586 761 587 771
rect 589 761 590 771
rect 629 761 630 771
rect 632 761 633 771
rect 1372 763 1373 773
rect 1375 763 1376 773
rect 1408 763 1409 773
rect 1411 763 1412 773
rect 1416 763 1417 773
rect 1419 763 1420 773
rect 1452 763 1453 773
rect 1455 763 1456 773
rect 1460 763 1461 773
rect 1463 763 1464 773
rect 1503 763 1504 773
rect 1506 763 1507 773
rect 1589 768 1590 778
rect 1592 768 1593 778
rect 743 719 744 732
rect 746 719 754 732
rect 756 719 757 732
rect 785 730 786 737
rect 788 730 789 737
rect 1176 717 1177 723
rect 1179 717 1180 723
rect 1003 685 1004 695
rect 1006 685 1007 695
rect 505 661 506 671
rect 508 661 509 671
rect 541 661 542 671
rect 544 661 545 671
rect 549 661 550 671
rect 552 661 553 671
rect 585 661 586 671
rect 588 661 589 671
rect 593 661 594 671
rect 596 661 597 671
rect 636 661 637 671
rect 639 661 640 671
rect 1215 668 1216 680
rect 1218 668 1226 680
rect 1228 668 1229 680
rect 1243 668 1244 680
rect 1246 668 1254 680
rect 1256 668 1257 680
rect 929 615 930 656
rect 932 615 937 656
rect 939 615 940 656
rect 962 616 963 656
rect 965 616 966 656
rect 989 616 990 656
rect 992 616 993 656
rect 1176 662 1177 668
rect 1179 662 1180 668
rect 1591 669 1592 679
rect 1594 669 1595 679
rect 1371 656 1372 666
rect 1374 656 1375 666
rect 1407 656 1408 666
rect 1410 656 1411 666
rect 1415 656 1416 666
rect 1418 656 1419 666
rect 1451 656 1452 666
rect 1454 656 1455 666
rect 1459 656 1460 666
rect 1462 656 1463 666
rect 1502 656 1503 666
rect 1505 656 1506 666
rect 516 547 517 557
rect 519 547 520 557
rect 552 547 553 557
rect 555 547 556 557
rect 560 547 561 557
rect 563 547 564 557
rect 596 547 597 557
rect 599 547 600 557
rect 604 547 605 557
rect 607 547 608 557
rect 647 547 648 557
rect 650 547 651 557
rect 915 538 916 578
rect 918 538 919 578
rect 939 538 940 578
rect 942 538 943 578
rect 960 538 961 578
rect 963 538 964 578
rect 977 538 978 578
rect 980 538 981 578
rect 1179 593 1180 599
rect 1182 593 1183 599
rect 1017 536 1018 546
rect 1020 536 1021 546
rect 1587 567 1588 577
rect 1590 567 1591 577
rect 1218 544 1219 556
rect 1221 544 1229 556
rect 1231 544 1232 556
rect 1246 544 1247 556
rect 1249 544 1257 556
rect 1259 544 1260 556
rect 1371 552 1372 562
rect 1374 552 1375 562
rect 1407 552 1408 562
rect 1410 552 1411 562
rect 1415 552 1416 562
rect 1418 552 1419 562
rect 1451 552 1452 562
rect 1454 552 1455 562
rect 1459 552 1460 562
rect 1462 552 1463 562
rect 1502 552 1503 562
rect 1505 552 1506 562
rect 1179 538 1180 544
rect 1182 538 1183 544
rect 1008 458 1009 468
rect 1011 458 1012 468
rect 508 438 509 448
rect 511 438 512 448
rect 544 438 545 448
rect 547 438 548 448
rect 552 438 553 448
rect 555 438 556 448
rect 588 438 589 448
rect 591 438 592 448
rect 596 438 597 448
rect 599 438 600 448
rect 639 438 640 448
rect 642 438 643 448
rect 1173 445 1174 451
rect 1176 445 1177 451
rect 961 388 962 429
rect 964 388 969 429
rect 971 388 972 429
rect 994 389 995 429
rect 997 389 998 429
rect 1584 448 1585 458
rect 1587 448 1588 458
rect 1371 437 1372 447
rect 1374 437 1375 447
rect 1407 437 1408 447
rect 1410 437 1411 447
rect 1415 437 1416 447
rect 1418 437 1419 447
rect 1451 437 1452 447
rect 1454 437 1455 447
rect 1459 437 1460 447
rect 1462 437 1463 447
rect 1502 437 1503 447
rect 1505 437 1506 447
rect 1212 396 1213 408
rect 1215 396 1223 408
rect 1225 396 1226 408
rect 1240 396 1241 408
rect 1243 396 1251 408
rect 1253 396 1254 408
rect 1173 390 1174 396
rect 1176 390 1177 396
rect 513 313 514 323
rect 516 313 517 323
rect 549 313 550 323
rect 552 313 553 323
rect 557 313 558 323
rect 560 313 561 323
rect 593 313 594 323
rect 596 313 597 323
rect 601 313 602 323
rect 604 313 605 323
rect 644 313 645 323
rect 647 313 648 323
rect 947 311 948 351
rect 950 311 951 351
rect 971 311 972 351
rect 974 311 975 351
rect 992 311 993 351
rect 995 311 996 351
rect 1022 309 1023 319
rect 1025 309 1026 319
rect 1010 235 1011 245
rect 1013 235 1014 245
rect 529 202 530 212
rect 532 202 533 212
rect 565 202 566 212
rect 568 202 569 212
rect 573 202 574 212
rect 576 202 577 212
rect 609 202 610 212
rect 612 202 613 212
rect 617 202 618 212
rect 620 202 621 212
rect 660 202 661 212
rect 663 202 664 212
rect 982 165 983 206
rect 985 165 990 206
rect 992 165 993 206
rect 519 84 520 94
rect 522 84 523 94
rect 555 84 556 94
rect 558 84 559 94
rect 563 84 564 94
rect 566 84 567 94
rect 599 84 600 94
rect 602 84 603 94
rect 607 84 608 94
rect 610 84 611 94
rect 650 84 651 94
rect 653 84 654 94
rect 968 88 969 128
rect 971 88 972 128
rect 992 88 993 128
rect 995 88 996 128
rect 1024 86 1025 96
rect 1027 86 1028 96
<< pdiffusion >>
rect 816 1097 817 1109
rect 819 1097 820 1109
rect 855 1081 856 1105
rect 858 1081 860 1105
rect 864 1081 866 1105
rect 868 1081 869 1105
rect 883 1075 884 1099
rect 886 1075 888 1099
rect 892 1075 894 1099
rect 896 1075 897 1099
rect 956 1097 957 1109
rect 959 1097 960 1109
rect 995 1081 996 1105
rect 998 1081 1000 1105
rect 1004 1081 1006 1105
rect 1008 1081 1009 1105
rect 816 1042 817 1054
rect 819 1042 820 1054
rect 1023 1075 1024 1099
rect 1026 1075 1028 1099
rect 1032 1075 1034 1099
rect 1036 1075 1037 1099
rect 1091 1097 1092 1109
rect 1094 1097 1095 1109
rect 1130 1081 1131 1105
rect 1133 1081 1135 1105
rect 1139 1081 1141 1105
rect 1143 1081 1144 1105
rect 956 1042 957 1054
rect 959 1042 960 1054
rect 1158 1075 1159 1099
rect 1161 1075 1163 1099
rect 1167 1075 1169 1099
rect 1171 1075 1172 1099
rect 1229 1096 1230 1108
rect 1232 1096 1233 1108
rect 1268 1080 1269 1104
rect 1271 1080 1273 1104
rect 1277 1080 1279 1104
rect 1281 1080 1282 1104
rect 1091 1042 1092 1054
rect 1094 1042 1095 1054
rect 1296 1074 1297 1098
rect 1299 1074 1301 1098
rect 1305 1074 1307 1098
rect 1309 1074 1310 1098
rect 1229 1041 1230 1053
rect 1232 1041 1233 1053
rect 493 989 494 1014
rect 496 989 497 1014
rect 501 989 502 1014
rect 504 989 505 1014
rect 531 989 532 1014
rect 534 989 535 1014
rect 575 989 576 1014
rect 578 989 579 1014
rect 620 989 621 1014
rect 623 989 624 1014
rect 743 972 744 984
rect 746 972 748 984
rect 752 972 754 984
rect 756 972 757 984
rect 785 972 786 984
rect 788 972 789 984
rect 1007 951 1008 971
rect 1010 951 1011 971
rect 1178 970 1179 982
rect 1181 970 1182 982
rect 1217 954 1218 978
rect 1220 954 1222 978
rect 1226 954 1228 978
rect 1230 954 1231 978
rect 1245 948 1246 972
rect 1248 948 1250 972
rect 1254 948 1256 972
rect 1258 948 1259 972
rect 497 891 498 916
rect 500 891 501 916
rect 505 891 506 916
rect 508 891 509 916
rect 535 891 536 916
rect 538 891 539 916
rect 579 891 580 916
rect 582 891 583 916
rect 624 891 625 916
rect 627 891 628 916
rect 1178 915 1179 927
rect 1181 915 1182 927
rect 743 898 744 910
rect 746 898 748 910
rect 752 898 754 910
rect 756 898 757 910
rect 785 898 786 910
rect 788 898 789 910
rect 1037 861 1038 901
rect 1040 861 1041 901
rect 1378 895 1379 920
rect 1381 895 1382 920
rect 1386 895 1387 920
rect 1389 895 1390 920
rect 1416 895 1417 920
rect 1419 895 1420 920
rect 1460 895 1461 920
rect 1463 895 1464 920
rect 1505 895 1506 920
rect 1508 895 1509 920
rect 1585 899 1586 919
rect 1588 899 1589 919
rect 743 829 744 841
rect 746 829 748 841
rect 752 829 754 841
rect 756 829 757 841
rect 785 829 786 841
rect 788 829 789 841
rect 1074 833 1075 843
rect 1077 833 1078 843
rect 502 793 503 818
rect 505 793 506 818
rect 510 793 511 818
rect 513 793 514 818
rect 540 793 541 818
rect 543 793 544 818
rect 584 793 585 818
rect 587 793 588 818
rect 629 793 630 818
rect 632 793 633 818
rect 1021 802 1022 822
rect 1024 802 1025 822
rect 1376 795 1377 820
rect 1379 795 1380 820
rect 1384 795 1385 820
rect 1387 795 1388 820
rect 1414 795 1415 820
rect 1417 795 1418 820
rect 1458 795 1459 820
rect 1461 795 1462 820
rect 1503 795 1504 820
rect 1506 795 1507 820
rect 1589 796 1590 816
rect 1592 796 1593 816
rect 743 755 744 767
rect 746 755 748 767
rect 752 755 754 767
rect 756 755 757 767
rect 785 755 786 767
rect 788 755 789 767
rect 1176 737 1177 749
rect 1179 737 1180 749
rect 509 693 510 718
rect 512 693 513 718
rect 517 693 518 718
rect 520 693 521 718
rect 547 693 548 718
rect 550 693 551 718
rect 591 693 592 718
rect 594 693 595 718
rect 636 693 637 718
rect 639 693 640 718
rect 1003 713 1004 733
rect 1006 713 1007 733
rect 1215 721 1216 745
rect 1218 721 1220 745
rect 1224 721 1226 745
rect 1228 721 1229 745
rect 1243 715 1244 739
rect 1246 715 1248 739
rect 1252 715 1254 739
rect 1256 715 1257 739
rect 1176 682 1177 694
rect 1179 682 1180 694
rect 1375 688 1376 713
rect 1378 688 1379 713
rect 1383 688 1384 713
rect 1386 688 1387 713
rect 1413 688 1414 713
rect 1416 688 1417 713
rect 1457 688 1458 713
rect 1460 688 1461 713
rect 1502 688 1503 713
rect 1505 688 1506 713
rect 1591 697 1592 717
rect 1594 697 1595 717
rect 1033 623 1034 663
rect 1036 623 1037 663
rect 1179 613 1180 625
rect 1182 613 1183 625
rect 520 579 521 604
rect 523 579 524 604
rect 528 579 529 604
rect 531 579 532 604
rect 558 579 559 604
rect 561 579 562 604
rect 602 579 603 604
rect 605 579 606 604
rect 647 579 648 604
rect 650 579 651 604
rect 1070 595 1071 605
rect 1073 595 1074 605
rect 1017 564 1018 584
rect 1020 564 1021 584
rect 1218 597 1219 621
rect 1221 597 1223 621
rect 1227 597 1229 621
rect 1231 597 1232 621
rect 1246 591 1247 615
rect 1249 591 1251 615
rect 1255 591 1257 615
rect 1259 591 1260 615
rect 1179 558 1180 570
rect 1182 558 1183 570
rect 1375 584 1376 609
rect 1378 584 1379 609
rect 1383 584 1384 609
rect 1386 584 1387 609
rect 1413 584 1414 609
rect 1416 584 1417 609
rect 1457 584 1458 609
rect 1460 584 1461 609
rect 1502 584 1503 609
rect 1505 584 1506 609
rect 1587 595 1588 615
rect 1590 595 1591 615
rect 512 470 513 495
rect 515 470 516 495
rect 520 470 521 495
rect 523 470 524 495
rect 550 470 551 495
rect 553 470 554 495
rect 594 470 595 495
rect 597 470 598 495
rect 639 470 640 495
rect 642 470 643 495
rect 1008 486 1009 506
rect 1011 486 1012 506
rect 1173 465 1174 477
rect 1176 465 1177 477
rect 1212 449 1213 473
rect 1215 449 1217 473
rect 1221 449 1223 473
rect 1225 449 1226 473
rect 1375 469 1376 494
rect 1378 469 1379 494
rect 1383 469 1384 494
rect 1386 469 1387 494
rect 1413 469 1414 494
rect 1416 469 1417 494
rect 1457 469 1458 494
rect 1460 469 1461 494
rect 1502 469 1503 494
rect 1505 469 1506 494
rect 1584 476 1585 496
rect 1587 476 1588 496
rect 1038 396 1039 436
rect 1041 396 1042 436
rect 1240 443 1241 467
rect 1243 443 1245 467
rect 1249 443 1251 467
rect 1253 443 1254 467
rect 1173 410 1174 422
rect 1176 410 1177 422
rect 517 345 518 370
rect 520 345 521 370
rect 525 345 526 370
rect 528 345 529 370
rect 555 345 556 370
rect 558 345 559 370
rect 599 345 600 370
rect 602 345 603 370
rect 644 345 645 370
rect 647 345 648 370
rect 1075 368 1076 378
rect 1078 368 1079 378
rect 1022 337 1023 357
rect 1025 337 1026 357
rect 1010 263 1011 283
rect 1013 263 1014 283
rect 533 234 534 259
rect 536 234 537 259
rect 541 234 542 259
rect 544 234 545 259
rect 571 234 572 259
rect 574 234 575 259
rect 615 234 616 259
rect 618 234 619 259
rect 660 234 661 259
rect 663 234 664 259
rect 1040 173 1041 213
rect 1043 173 1044 213
rect 1077 145 1078 155
rect 1080 145 1081 155
rect 523 116 524 141
rect 526 116 527 141
rect 531 116 532 141
rect 534 116 535 141
rect 561 116 562 141
rect 564 116 565 141
rect 605 116 606 141
rect 608 116 609 141
rect 650 116 651 141
rect 653 116 654 141
rect 1024 114 1025 134
rect 1027 114 1028 134
<< ndcontact >>
rect 812 1077 816 1083
rect 820 1077 824 1083
rect 952 1077 956 1083
rect 960 1077 964 1083
rect 1087 1077 1091 1083
rect 1095 1077 1099 1083
rect 851 1028 855 1040
rect 869 1028 873 1040
rect 879 1028 883 1040
rect 897 1028 901 1040
rect 1225 1076 1229 1082
rect 1233 1076 1237 1082
rect 991 1028 995 1040
rect 1009 1028 1013 1040
rect 1019 1028 1023 1040
rect 1037 1028 1041 1040
rect 1126 1028 1130 1040
rect 1144 1028 1148 1040
rect 1154 1028 1158 1040
rect 1172 1028 1176 1040
rect 812 1022 816 1028
rect 820 1022 824 1028
rect 952 1022 956 1028
rect 960 1022 964 1028
rect 1087 1022 1091 1028
rect 1095 1022 1099 1028
rect 1264 1027 1268 1039
rect 1282 1027 1286 1039
rect 1292 1027 1296 1039
rect 1310 1027 1314 1039
rect 1225 1021 1229 1027
rect 1233 1021 1237 1027
rect 485 957 489 967
rect 493 957 497 967
rect 521 957 525 967
rect 529 957 533 967
rect 537 957 541 967
rect 565 957 569 967
rect 573 957 577 967
rect 581 957 585 967
rect 616 957 620 967
rect 624 957 628 967
rect 739 936 743 949
rect 757 936 761 949
rect 781 947 785 954
rect 789 947 793 954
rect 1174 950 1178 956
rect 1182 950 1186 956
rect 1003 923 1007 933
rect 1011 923 1015 933
rect 1213 901 1217 913
rect 1231 901 1235 913
rect 1241 901 1245 913
rect 1259 901 1263 913
rect 489 859 493 869
rect 497 859 501 869
rect 525 859 529 869
rect 533 859 537 869
rect 541 859 545 869
rect 569 859 573 869
rect 577 859 581 869
rect 585 859 589 869
rect 620 859 624 869
rect 628 859 632 869
rect 739 862 743 875
rect 757 862 761 875
rect 781 873 785 880
rect 789 873 793 880
rect 912 853 916 894
rect 927 853 932 894
rect 945 854 949 894
rect 953 854 957 894
rect 972 854 976 894
rect 980 854 984 894
rect 995 854 999 894
rect 1003 854 1007 894
rect 1174 895 1178 901
rect 1182 895 1186 901
rect 1370 863 1374 873
rect 1378 863 1382 873
rect 1406 863 1410 873
rect 1414 863 1418 873
rect 1422 863 1426 873
rect 1450 863 1454 873
rect 1458 863 1462 873
rect 1466 863 1470 873
rect 1501 863 1505 873
rect 1509 863 1513 873
rect 1581 871 1585 881
rect 1589 871 1593 881
rect 739 793 743 806
rect 757 793 761 806
rect 781 804 785 811
rect 789 804 793 811
rect 898 776 902 816
rect 906 776 910 816
rect 922 776 926 816
rect 930 776 934 816
rect 943 776 947 816
rect 951 776 955 816
rect 960 776 964 816
rect 968 776 972 816
rect 978 777 982 817
rect 986 777 990 817
rect 1017 774 1021 784
rect 1025 774 1029 784
rect 494 761 498 771
rect 502 761 506 771
rect 530 761 534 771
rect 538 761 542 771
rect 546 761 550 771
rect 574 761 578 771
rect 582 761 586 771
rect 590 761 594 771
rect 625 761 629 771
rect 633 761 637 771
rect 1368 763 1372 773
rect 1376 763 1380 773
rect 1404 763 1408 773
rect 1412 763 1416 773
rect 1420 763 1424 773
rect 1448 763 1452 773
rect 1456 763 1460 773
rect 1464 763 1468 773
rect 1499 763 1503 773
rect 1507 763 1511 773
rect 1585 768 1589 778
rect 1593 768 1597 778
rect 739 719 743 732
rect 757 719 761 732
rect 781 730 785 737
rect 789 730 793 737
rect 1172 717 1176 723
rect 1180 717 1184 723
rect 999 685 1003 695
rect 1007 685 1011 695
rect 501 661 505 671
rect 509 661 513 671
rect 537 661 541 671
rect 545 661 549 671
rect 553 661 557 671
rect 581 661 585 671
rect 589 661 593 671
rect 597 661 601 671
rect 632 661 636 671
rect 640 661 644 671
rect 1211 668 1215 680
rect 1229 668 1233 680
rect 1239 668 1243 680
rect 1257 668 1261 680
rect 925 615 929 656
rect 940 615 945 656
rect 958 616 962 656
rect 966 616 970 656
rect 985 616 989 656
rect 993 616 997 656
rect 1172 662 1176 668
rect 1180 662 1184 668
rect 1587 669 1591 679
rect 1595 669 1599 679
rect 1367 656 1371 666
rect 1375 656 1379 666
rect 1403 656 1407 666
rect 1411 656 1415 666
rect 1419 656 1423 666
rect 1447 656 1451 666
rect 1455 656 1459 666
rect 1463 656 1467 666
rect 1498 656 1502 666
rect 1506 656 1510 666
rect 512 547 516 557
rect 520 547 524 557
rect 548 547 552 557
rect 556 547 560 557
rect 564 547 568 557
rect 592 547 596 557
rect 600 547 604 557
rect 608 547 612 557
rect 643 547 647 557
rect 651 547 655 557
rect 911 538 915 578
rect 919 538 923 578
rect 935 538 939 578
rect 943 538 947 578
rect 956 538 960 578
rect 964 538 968 578
rect 973 538 977 578
rect 981 538 985 578
rect 1175 593 1179 599
rect 1183 593 1187 599
rect 1013 536 1017 546
rect 1021 536 1025 546
rect 1583 567 1587 577
rect 1591 567 1595 577
rect 1214 544 1218 556
rect 1232 544 1236 556
rect 1242 544 1246 556
rect 1260 544 1264 556
rect 1367 552 1371 562
rect 1375 552 1379 562
rect 1403 552 1407 562
rect 1411 552 1415 562
rect 1419 552 1423 562
rect 1447 552 1451 562
rect 1455 552 1459 562
rect 1463 552 1467 562
rect 1498 552 1502 562
rect 1506 552 1510 562
rect 1175 538 1179 544
rect 1183 538 1187 544
rect 1004 458 1008 468
rect 1012 458 1016 468
rect 504 438 508 448
rect 512 438 516 448
rect 540 438 544 448
rect 548 438 552 448
rect 556 438 560 448
rect 584 438 588 448
rect 592 438 596 448
rect 600 438 604 448
rect 635 438 639 448
rect 643 438 647 448
rect 1169 445 1173 451
rect 1177 445 1181 451
rect 957 388 961 429
rect 972 388 977 429
rect 990 389 994 429
rect 998 389 1002 429
rect 1580 448 1584 458
rect 1588 448 1592 458
rect 1367 437 1371 447
rect 1375 437 1379 447
rect 1403 437 1407 447
rect 1411 437 1415 447
rect 1419 437 1423 447
rect 1447 437 1451 447
rect 1455 437 1459 447
rect 1463 437 1467 447
rect 1498 437 1502 447
rect 1506 437 1510 447
rect 1208 396 1212 408
rect 1226 396 1230 408
rect 1236 396 1240 408
rect 1254 396 1258 408
rect 1169 390 1173 396
rect 1177 390 1181 396
rect 509 313 513 323
rect 517 313 521 323
rect 545 313 549 323
rect 553 313 557 323
rect 561 313 565 323
rect 589 313 593 323
rect 597 313 601 323
rect 605 313 609 323
rect 640 313 644 323
rect 648 313 652 323
rect 943 311 947 351
rect 951 311 955 351
rect 967 311 971 351
rect 975 311 979 351
rect 988 311 992 351
rect 996 311 1000 351
rect 1018 309 1022 319
rect 1026 309 1030 319
rect 1006 235 1010 245
rect 1014 235 1018 245
rect 525 202 529 212
rect 533 202 537 212
rect 561 202 565 212
rect 569 202 573 212
rect 577 202 581 212
rect 605 202 609 212
rect 613 202 617 212
rect 621 202 625 212
rect 656 202 660 212
rect 664 202 668 212
rect 978 165 982 206
rect 993 165 998 206
rect 515 84 519 94
rect 523 84 527 94
rect 551 84 555 94
rect 559 84 563 94
rect 567 84 571 94
rect 595 84 599 94
rect 603 84 607 94
rect 611 84 615 94
rect 646 84 650 94
rect 654 84 658 94
rect 964 88 968 128
rect 972 88 976 128
rect 988 88 992 128
rect 996 88 1000 128
rect 1020 86 1024 96
rect 1028 86 1032 96
<< pdcontact >>
rect 812 1097 816 1109
rect 820 1097 824 1109
rect 851 1081 855 1105
rect 860 1081 864 1105
rect 869 1081 873 1105
rect 879 1075 883 1099
rect 888 1075 892 1099
rect 897 1075 901 1099
rect 952 1097 956 1109
rect 960 1097 964 1109
rect 991 1081 995 1105
rect 1000 1081 1004 1105
rect 1009 1081 1013 1105
rect 812 1042 816 1054
rect 820 1042 824 1054
rect 1019 1075 1023 1099
rect 1028 1075 1032 1099
rect 1037 1075 1041 1099
rect 1087 1097 1091 1109
rect 1095 1097 1099 1109
rect 1126 1081 1130 1105
rect 1135 1081 1139 1105
rect 1144 1081 1148 1105
rect 952 1042 956 1054
rect 960 1042 964 1054
rect 1154 1075 1158 1099
rect 1163 1075 1167 1099
rect 1172 1075 1176 1099
rect 1225 1096 1229 1108
rect 1233 1096 1237 1108
rect 1264 1080 1268 1104
rect 1273 1080 1277 1104
rect 1282 1080 1286 1104
rect 1087 1042 1091 1054
rect 1095 1042 1099 1054
rect 1292 1074 1296 1098
rect 1301 1074 1305 1098
rect 1310 1074 1314 1098
rect 1225 1041 1229 1053
rect 1233 1041 1237 1053
rect 489 989 493 1014
rect 497 989 501 1014
rect 505 989 509 1014
rect 527 989 531 1014
rect 535 989 539 1014
rect 571 989 575 1014
rect 579 989 583 1014
rect 616 989 620 1014
rect 624 989 628 1014
rect 739 972 743 984
rect 748 972 752 984
rect 757 972 761 984
rect 781 972 785 984
rect 789 972 793 984
rect 1003 951 1007 971
rect 1011 951 1015 971
rect 1174 970 1178 982
rect 1182 970 1186 982
rect 1213 954 1217 978
rect 1222 954 1226 978
rect 1231 954 1235 978
rect 1241 948 1245 972
rect 1250 948 1254 972
rect 1259 948 1263 972
rect 493 891 497 916
rect 501 891 505 916
rect 509 891 513 916
rect 531 891 535 916
rect 539 891 543 916
rect 575 891 579 916
rect 583 891 587 916
rect 620 891 624 916
rect 628 891 632 916
rect 1174 915 1178 927
rect 1182 915 1186 927
rect 739 898 743 910
rect 748 898 752 910
rect 757 898 761 910
rect 781 898 785 910
rect 789 898 793 910
rect 1033 861 1037 901
rect 1041 861 1045 901
rect 1374 895 1378 920
rect 1382 895 1386 920
rect 1390 895 1394 920
rect 1412 895 1416 920
rect 1420 895 1424 920
rect 1456 895 1460 920
rect 1464 895 1468 920
rect 1501 895 1505 920
rect 1509 895 1513 920
rect 1581 899 1585 919
rect 1589 899 1593 919
rect 739 829 743 841
rect 748 829 752 841
rect 757 829 761 841
rect 781 829 785 841
rect 789 829 793 841
rect 1070 833 1074 843
rect 1078 833 1082 843
rect 498 793 502 818
rect 506 793 510 818
rect 514 793 518 818
rect 536 793 540 818
rect 544 793 548 818
rect 580 793 584 818
rect 588 793 592 818
rect 625 793 629 818
rect 633 793 637 818
rect 1017 802 1021 822
rect 1025 802 1029 822
rect 1372 795 1376 820
rect 1380 795 1384 820
rect 1388 795 1392 820
rect 1410 795 1414 820
rect 1418 795 1422 820
rect 1454 795 1458 820
rect 1462 795 1466 820
rect 1499 795 1503 820
rect 1507 795 1511 820
rect 1585 796 1589 816
rect 1593 796 1597 816
rect 739 755 743 767
rect 748 755 752 767
rect 757 755 761 767
rect 781 755 785 767
rect 789 755 793 767
rect 1172 737 1176 749
rect 1180 737 1184 749
rect 505 693 509 718
rect 513 693 517 718
rect 521 693 525 718
rect 543 693 547 718
rect 551 693 555 718
rect 587 693 591 718
rect 595 693 599 718
rect 632 693 636 718
rect 640 693 644 718
rect 999 713 1003 733
rect 1007 713 1011 733
rect 1211 721 1215 745
rect 1220 721 1224 745
rect 1229 721 1233 745
rect 1239 715 1243 739
rect 1248 715 1252 739
rect 1257 715 1261 739
rect 1172 682 1176 694
rect 1180 682 1184 694
rect 1371 688 1375 713
rect 1379 688 1383 713
rect 1387 688 1391 713
rect 1409 688 1413 713
rect 1417 688 1421 713
rect 1453 688 1457 713
rect 1461 688 1465 713
rect 1498 688 1502 713
rect 1506 688 1510 713
rect 1587 697 1591 717
rect 1595 697 1599 717
rect 1029 623 1033 663
rect 1037 623 1041 663
rect 1175 613 1179 625
rect 1183 613 1187 625
rect 516 579 520 604
rect 524 579 528 604
rect 532 579 536 604
rect 554 579 558 604
rect 562 579 566 604
rect 598 579 602 604
rect 606 579 610 604
rect 643 579 647 604
rect 651 579 655 604
rect 1066 595 1070 605
rect 1074 595 1078 605
rect 1013 564 1017 584
rect 1021 564 1025 584
rect 1214 597 1218 621
rect 1223 597 1227 621
rect 1232 597 1236 621
rect 1242 591 1246 615
rect 1251 591 1255 615
rect 1260 591 1264 615
rect 1175 558 1179 570
rect 1183 558 1187 570
rect 1371 584 1375 609
rect 1379 584 1383 609
rect 1387 584 1391 609
rect 1409 584 1413 609
rect 1417 584 1421 609
rect 1453 584 1457 609
rect 1461 584 1465 609
rect 1498 584 1502 609
rect 1506 584 1510 609
rect 1583 595 1587 615
rect 1591 595 1595 615
rect 508 470 512 495
rect 516 470 520 495
rect 524 470 528 495
rect 546 470 550 495
rect 554 470 558 495
rect 590 470 594 495
rect 598 470 602 495
rect 635 470 639 495
rect 643 470 647 495
rect 1004 486 1008 506
rect 1012 486 1016 506
rect 1169 465 1173 477
rect 1177 465 1181 477
rect 1208 449 1212 473
rect 1217 449 1221 473
rect 1226 449 1230 473
rect 1371 469 1375 494
rect 1379 469 1383 494
rect 1387 469 1391 494
rect 1409 469 1413 494
rect 1417 469 1421 494
rect 1453 469 1457 494
rect 1461 469 1465 494
rect 1498 469 1502 494
rect 1506 469 1510 494
rect 1580 476 1584 496
rect 1588 476 1592 496
rect 1034 396 1038 436
rect 1042 396 1046 436
rect 1236 443 1240 467
rect 1245 443 1249 467
rect 1254 443 1258 467
rect 1169 410 1173 422
rect 1177 410 1181 422
rect 513 345 517 370
rect 521 345 525 370
rect 529 345 533 370
rect 551 345 555 370
rect 559 345 563 370
rect 595 345 599 370
rect 603 345 607 370
rect 640 345 644 370
rect 648 345 652 370
rect 1071 368 1075 378
rect 1079 368 1083 378
rect 1018 337 1022 357
rect 1026 337 1030 357
rect 1006 263 1010 283
rect 1014 263 1018 283
rect 529 234 533 259
rect 537 234 541 259
rect 545 234 549 259
rect 567 234 571 259
rect 575 234 579 259
rect 611 234 615 259
rect 619 234 623 259
rect 656 234 660 259
rect 664 234 668 259
rect 1036 173 1040 213
rect 1044 173 1048 213
rect 1073 145 1077 155
rect 1081 145 1085 155
rect 519 116 523 141
rect 527 116 531 141
rect 535 116 539 141
rect 557 116 561 141
rect 565 116 569 141
rect 601 116 605 141
rect 609 116 613 141
rect 646 116 650 141
rect 654 116 658 141
rect 1020 114 1024 134
rect 1028 114 1032 134
<< polysilicon >>
rect 817 1109 819 1112
rect 957 1109 959 1112
rect 1092 1109 1094 1112
rect 856 1105 858 1108
rect 866 1105 868 1108
rect 817 1083 819 1097
rect 884 1099 886 1102
rect 894 1099 896 1102
rect 817 1074 819 1077
rect 856 1072 858 1081
rect 866 1071 868 1081
rect 996 1105 998 1108
rect 1006 1105 1008 1108
rect 957 1083 959 1097
rect 1024 1099 1026 1102
rect 1034 1099 1036 1102
rect 817 1054 819 1057
rect 817 1028 819 1042
rect 856 1040 858 1067
rect 866 1040 868 1066
rect 884 1064 886 1075
rect 884 1040 886 1060
rect 894 1053 896 1075
rect 957 1074 959 1077
rect 996 1072 998 1081
rect 1006 1071 1008 1081
rect 1230 1108 1232 1111
rect 1131 1105 1133 1108
rect 1141 1105 1143 1108
rect 1092 1083 1094 1097
rect 1159 1099 1161 1102
rect 1169 1099 1171 1102
rect 957 1054 959 1057
rect 894 1040 896 1049
rect 957 1028 959 1042
rect 996 1040 998 1067
rect 1006 1040 1008 1066
rect 1024 1064 1026 1075
rect 1024 1040 1026 1060
rect 1034 1053 1036 1075
rect 1092 1074 1094 1077
rect 1131 1072 1133 1081
rect 1141 1071 1143 1081
rect 1269 1104 1271 1107
rect 1279 1104 1281 1107
rect 1230 1082 1232 1096
rect 1297 1098 1299 1101
rect 1307 1098 1309 1101
rect 1092 1054 1094 1057
rect 1034 1040 1036 1049
rect 1092 1028 1094 1042
rect 1131 1040 1133 1067
rect 1141 1040 1143 1066
rect 1159 1064 1161 1075
rect 1159 1040 1161 1060
rect 1169 1053 1171 1075
rect 1230 1073 1232 1076
rect 1269 1071 1271 1080
rect 1279 1070 1281 1080
rect 1230 1053 1232 1056
rect 1169 1040 1171 1049
rect 856 1025 858 1028
rect 866 1025 868 1028
rect 884 1025 886 1028
rect 894 1025 896 1028
rect 996 1025 998 1028
rect 1006 1025 1008 1028
rect 1024 1025 1026 1028
rect 1034 1025 1036 1028
rect 1131 1025 1133 1028
rect 1141 1025 1143 1028
rect 1159 1025 1161 1028
rect 1169 1025 1171 1028
rect 1230 1027 1232 1041
rect 1269 1039 1271 1066
rect 1279 1039 1281 1065
rect 1297 1063 1299 1074
rect 1297 1039 1299 1059
rect 1307 1052 1309 1074
rect 1307 1039 1309 1048
rect 817 1019 819 1022
rect 957 1019 959 1022
rect 1092 1019 1094 1022
rect 1269 1024 1271 1027
rect 1279 1024 1281 1027
rect 1297 1024 1299 1027
rect 1307 1024 1309 1027
rect 1230 1018 1232 1021
rect 494 1014 496 1017
rect 502 1014 504 1017
rect 532 1014 534 1017
rect 576 1014 578 1017
rect 621 1014 623 1017
rect 494 982 496 989
rect 489 978 496 982
rect 490 967 492 978
rect 502 970 504 989
rect 532 981 534 989
rect 576 981 578 989
rect 526 979 534 981
rect 570 979 578 981
rect 526 967 528 979
rect 534 967 536 976
rect 570 967 572 979
rect 578 967 580 976
rect 621 967 623 989
rect 744 984 746 987
rect 754 984 756 987
rect 786 984 788 987
rect 1179 982 1181 985
rect 490 954 492 957
rect 526 954 528 957
rect 534 954 536 957
rect 570 954 572 957
rect 578 954 580 957
rect 621 954 623 957
rect 744 949 746 972
rect 754 949 756 972
rect 786 954 788 972
rect 1008 971 1010 974
rect 1218 978 1220 981
rect 1228 978 1230 981
rect 1179 956 1181 970
rect 786 944 788 947
rect 744 932 746 936
rect 754 932 756 936
rect 1008 933 1010 951
rect 1246 972 1248 975
rect 1256 972 1258 975
rect 1179 947 1181 950
rect 1218 945 1220 954
rect 1228 944 1230 954
rect 1179 927 1181 930
rect 1008 920 1010 923
rect 498 916 500 919
rect 506 916 508 919
rect 536 916 538 919
rect 580 916 582 919
rect 625 916 627 919
rect 744 910 746 913
rect 754 910 756 913
rect 786 910 788 913
rect 1038 901 1040 904
rect 1179 901 1181 915
rect 1218 913 1220 940
rect 1228 913 1230 939
rect 1246 937 1248 948
rect 1246 913 1248 933
rect 1256 926 1258 948
rect 1256 913 1258 922
rect 1379 920 1381 923
rect 1387 920 1389 923
rect 1417 920 1419 923
rect 1461 920 1463 923
rect 1506 920 1508 923
rect 498 884 500 891
rect 493 880 500 884
rect 494 869 496 880
rect 506 872 508 891
rect 536 883 538 891
rect 580 883 582 891
rect 530 881 538 883
rect 574 881 582 883
rect 530 869 532 881
rect 538 869 540 878
rect 574 869 576 881
rect 582 869 584 878
rect 625 869 627 891
rect 744 875 746 898
rect 754 875 756 898
rect 786 880 788 898
rect 917 894 919 901
rect 924 894 926 901
rect 950 894 952 901
rect 977 894 979 901
rect 1000 894 1002 901
rect 786 870 788 873
rect 494 856 496 859
rect 530 856 532 859
rect 538 856 540 859
rect 574 856 576 859
rect 582 856 584 859
rect 625 856 627 859
rect 744 858 746 862
rect 754 858 756 862
rect 1218 898 1220 901
rect 1228 898 1230 901
rect 1246 898 1248 901
rect 1256 898 1258 901
rect 1586 919 1588 922
rect 1179 892 1181 895
rect 1379 888 1381 895
rect 1374 884 1381 888
rect 1375 873 1377 884
rect 1387 876 1389 895
rect 1417 887 1419 895
rect 1461 887 1463 895
rect 1411 885 1419 887
rect 1455 885 1463 887
rect 1411 873 1413 885
rect 1419 873 1421 882
rect 1455 873 1457 885
rect 1463 873 1465 882
rect 1506 873 1508 895
rect 1586 881 1588 899
rect 1586 868 1588 871
rect 917 850 919 853
rect 924 850 926 853
rect 950 850 952 854
rect 977 850 979 854
rect 1000 850 1002 854
rect 1038 846 1040 861
rect 1375 860 1377 863
rect 1411 860 1413 863
rect 1419 860 1421 863
rect 1455 860 1457 863
rect 1463 860 1465 863
rect 1506 860 1508 863
rect 744 841 746 844
rect 754 841 756 844
rect 786 841 788 844
rect 1075 843 1077 846
rect 503 818 505 821
rect 511 818 513 821
rect 541 818 543 821
rect 585 818 587 821
rect 630 818 632 821
rect 744 806 746 829
rect 754 806 756 829
rect 786 811 788 829
rect 903 816 905 823
rect 927 816 929 823
rect 948 816 950 823
rect 965 816 967 823
rect 983 817 985 824
rect 1022 822 1024 825
rect 786 801 788 804
rect 503 786 505 793
rect 498 782 505 786
rect 499 771 501 782
rect 511 774 513 793
rect 541 785 543 793
rect 585 785 587 793
rect 535 783 543 785
rect 579 783 587 785
rect 535 771 537 783
rect 543 771 545 780
rect 579 771 581 783
rect 587 771 589 780
rect 630 771 632 793
rect 744 789 746 793
rect 754 789 756 793
rect 1075 818 1077 833
rect 1377 820 1379 823
rect 1385 820 1387 823
rect 1415 820 1417 823
rect 1459 820 1461 823
rect 1504 820 1506 823
rect 1022 784 1024 802
rect 1590 816 1592 819
rect 1377 788 1379 795
rect 1372 784 1379 788
rect 903 772 905 776
rect 927 772 929 776
rect 948 772 950 776
rect 965 772 967 776
rect 983 773 985 777
rect 1022 771 1024 774
rect 1373 773 1375 784
rect 1385 776 1387 795
rect 1415 787 1417 795
rect 1459 787 1461 795
rect 1409 785 1417 787
rect 1453 785 1461 787
rect 1409 773 1411 785
rect 1417 773 1419 782
rect 1453 773 1455 785
rect 1461 773 1463 782
rect 1504 773 1506 795
rect 1590 778 1592 796
rect 744 767 746 770
rect 754 767 756 770
rect 786 767 788 770
rect 499 758 501 761
rect 535 758 537 761
rect 543 758 545 761
rect 579 758 581 761
rect 587 758 589 761
rect 630 758 632 761
rect 1590 765 1592 768
rect 1373 760 1375 763
rect 1409 760 1411 763
rect 1417 760 1419 763
rect 1453 760 1455 763
rect 1461 760 1463 763
rect 1504 760 1506 763
rect 744 732 746 755
rect 754 732 756 755
rect 786 737 788 755
rect 1177 749 1179 752
rect 1216 745 1218 748
rect 1226 745 1228 748
rect 510 718 512 721
rect 518 718 520 721
rect 548 718 550 721
rect 592 718 594 721
rect 637 718 639 721
rect 1004 733 1006 736
rect 786 727 788 730
rect 744 715 746 719
rect 754 715 756 719
rect 1177 723 1179 737
rect 1244 739 1246 742
rect 1254 739 1256 742
rect 1177 714 1179 717
rect 1004 695 1006 713
rect 1216 712 1218 721
rect 1226 711 1228 721
rect 1592 717 1594 720
rect 510 686 512 693
rect 505 682 512 686
rect 506 671 508 682
rect 518 674 520 693
rect 548 685 550 693
rect 592 685 594 693
rect 542 683 550 685
rect 586 683 594 685
rect 542 671 544 683
rect 550 671 552 680
rect 586 671 588 683
rect 594 671 596 680
rect 637 671 639 693
rect 1177 694 1179 697
rect 1004 682 1006 685
rect 1177 668 1179 682
rect 1216 680 1218 707
rect 1226 680 1228 706
rect 1244 704 1246 715
rect 1244 680 1246 700
rect 1254 693 1256 715
rect 1376 713 1378 716
rect 1384 713 1386 716
rect 1414 713 1416 716
rect 1458 713 1460 716
rect 1503 713 1505 716
rect 1254 680 1256 689
rect 1376 681 1378 688
rect 1371 677 1378 681
rect 1034 663 1036 666
rect 506 658 508 661
rect 542 658 544 661
rect 550 658 552 661
rect 586 658 588 661
rect 594 658 596 661
rect 637 658 639 661
rect 930 656 932 663
rect 937 656 939 663
rect 963 656 965 663
rect 990 656 992 663
rect 1216 665 1218 668
rect 1226 665 1228 668
rect 1244 665 1246 668
rect 1254 665 1256 668
rect 1372 666 1374 677
rect 1384 669 1386 688
rect 1414 680 1416 688
rect 1458 680 1460 688
rect 1408 678 1416 680
rect 1452 678 1460 680
rect 1408 666 1410 678
rect 1416 666 1418 675
rect 1452 666 1454 678
rect 1460 666 1462 675
rect 1503 666 1505 688
rect 1592 679 1594 697
rect 1592 666 1594 669
rect 1177 659 1179 662
rect 1372 653 1374 656
rect 1408 653 1410 656
rect 1416 653 1418 656
rect 1452 653 1454 656
rect 1460 653 1462 656
rect 1503 653 1505 656
rect 1180 625 1182 628
rect 930 612 932 615
rect 937 612 939 615
rect 963 612 965 616
rect 990 612 992 616
rect 1034 608 1036 623
rect 1219 621 1221 624
rect 1229 621 1231 624
rect 521 604 523 607
rect 529 604 531 607
rect 559 604 561 607
rect 603 604 605 607
rect 648 604 650 607
rect 1071 605 1073 608
rect 1180 599 1182 613
rect 521 572 523 579
rect 516 568 523 572
rect 517 557 519 568
rect 529 560 531 579
rect 559 571 561 579
rect 603 571 605 579
rect 553 569 561 571
rect 597 569 605 571
rect 553 557 555 569
rect 561 557 563 566
rect 597 557 599 569
rect 605 557 607 566
rect 648 557 650 579
rect 916 578 918 585
rect 940 578 942 585
rect 961 578 963 585
rect 978 578 980 585
rect 1018 584 1020 587
rect 517 544 519 547
rect 553 544 555 547
rect 561 544 563 547
rect 597 544 599 547
rect 605 544 607 547
rect 648 544 650 547
rect 1071 580 1073 595
rect 1247 615 1249 618
rect 1257 615 1259 618
rect 1588 615 1590 618
rect 1180 590 1182 593
rect 1219 588 1221 597
rect 1229 587 1231 597
rect 1376 609 1378 612
rect 1384 609 1386 612
rect 1414 609 1416 612
rect 1458 609 1460 612
rect 1503 609 1505 612
rect 1180 570 1182 573
rect 1018 546 1020 564
rect 916 534 918 538
rect 940 534 942 538
rect 961 534 963 538
rect 978 534 980 538
rect 1180 544 1182 558
rect 1219 556 1221 583
rect 1229 556 1231 582
rect 1247 580 1249 591
rect 1247 556 1249 576
rect 1257 569 1259 591
rect 1376 577 1378 584
rect 1371 573 1378 577
rect 1257 556 1259 565
rect 1372 562 1374 573
rect 1384 565 1386 584
rect 1414 576 1416 584
rect 1458 576 1460 584
rect 1408 574 1416 576
rect 1452 574 1460 576
rect 1408 562 1410 574
rect 1416 562 1418 571
rect 1452 562 1454 574
rect 1460 562 1462 571
rect 1503 562 1505 584
rect 1588 577 1590 595
rect 1588 564 1590 567
rect 1372 549 1374 552
rect 1408 549 1410 552
rect 1416 549 1418 552
rect 1452 549 1454 552
rect 1460 549 1462 552
rect 1503 549 1505 552
rect 1219 541 1221 544
rect 1229 541 1231 544
rect 1247 541 1249 544
rect 1257 541 1259 544
rect 1018 533 1020 536
rect 1180 535 1182 538
rect 1009 506 1011 509
rect 513 495 515 498
rect 521 495 523 498
rect 551 495 553 498
rect 595 495 597 498
rect 640 495 642 498
rect 1376 494 1378 497
rect 1384 494 1386 497
rect 1414 494 1416 497
rect 1458 494 1460 497
rect 1503 494 1505 497
rect 1585 496 1587 499
rect 513 463 515 470
rect 508 459 515 463
rect 509 448 511 459
rect 521 451 523 470
rect 551 462 553 470
rect 595 462 597 470
rect 545 460 553 462
rect 589 460 597 462
rect 545 448 547 460
rect 553 448 555 457
rect 589 448 591 460
rect 597 448 599 457
rect 640 448 642 470
rect 1009 468 1011 486
rect 1174 477 1176 480
rect 1213 473 1215 476
rect 1223 473 1225 476
rect 1009 455 1011 458
rect 1174 451 1176 465
rect 1241 467 1243 470
rect 1251 467 1253 470
rect 1174 442 1176 445
rect 1213 440 1215 449
rect 509 435 511 438
rect 545 435 547 438
rect 553 435 555 438
rect 589 435 591 438
rect 597 435 599 438
rect 640 435 642 438
rect 1039 436 1041 439
rect 962 429 964 436
rect 969 429 971 436
rect 995 429 997 436
rect 1223 439 1225 449
rect 1376 462 1378 469
rect 1371 458 1378 462
rect 1372 447 1374 458
rect 1384 450 1386 469
rect 1414 461 1416 469
rect 1458 461 1460 469
rect 1408 459 1416 461
rect 1452 459 1460 461
rect 1408 447 1410 459
rect 1416 447 1418 456
rect 1452 447 1454 459
rect 1460 447 1462 456
rect 1503 447 1505 469
rect 1585 458 1587 476
rect 1174 422 1176 425
rect 1174 396 1176 410
rect 1213 408 1215 435
rect 1223 408 1225 434
rect 1241 432 1243 443
rect 1241 408 1243 428
rect 1251 421 1253 443
rect 1585 445 1587 448
rect 1372 434 1374 437
rect 1408 434 1410 437
rect 1416 434 1418 437
rect 1452 434 1454 437
rect 1460 434 1462 437
rect 1503 434 1505 437
rect 1251 408 1253 417
rect 962 385 964 388
rect 969 385 971 388
rect 995 385 997 389
rect 1039 381 1041 396
rect 1213 393 1215 396
rect 1223 393 1225 396
rect 1241 393 1243 396
rect 1251 393 1253 396
rect 1174 387 1176 390
rect 1076 378 1078 381
rect 518 370 520 373
rect 526 370 528 373
rect 556 370 558 373
rect 600 370 602 373
rect 645 370 647 373
rect 948 351 950 358
rect 972 351 974 358
rect 993 351 995 358
rect 1023 357 1025 360
rect 518 338 520 345
rect 513 334 520 338
rect 514 323 516 334
rect 526 326 528 345
rect 556 337 558 345
rect 600 337 602 345
rect 550 335 558 337
rect 594 335 602 337
rect 550 323 552 335
rect 558 323 560 332
rect 594 323 596 335
rect 602 323 604 332
rect 645 323 647 345
rect 514 310 516 313
rect 550 310 552 313
rect 558 310 560 313
rect 594 310 596 313
rect 602 310 604 313
rect 645 310 647 313
rect 1076 353 1078 368
rect 1023 319 1025 337
rect 948 307 950 311
rect 972 307 974 311
rect 993 307 995 311
rect 1023 306 1025 309
rect 1011 283 1013 286
rect 534 259 536 262
rect 542 259 544 262
rect 572 259 574 262
rect 616 259 618 262
rect 661 259 663 262
rect 1011 245 1013 263
rect 534 227 536 234
rect 529 223 536 227
rect 530 212 532 223
rect 542 215 544 234
rect 572 226 574 234
rect 616 226 618 234
rect 566 224 574 226
rect 610 224 618 226
rect 566 212 568 224
rect 574 212 576 221
rect 610 212 612 224
rect 618 212 620 221
rect 661 212 663 234
rect 1011 232 1013 235
rect 1041 213 1043 216
rect 983 206 985 213
rect 990 206 992 213
rect 530 199 532 202
rect 566 199 568 202
rect 574 199 576 202
rect 610 199 612 202
rect 618 199 620 202
rect 661 199 663 202
rect 983 162 985 165
rect 990 162 992 165
rect 1041 158 1043 173
rect 1078 155 1080 158
rect 524 141 526 144
rect 532 141 534 144
rect 562 141 564 144
rect 606 141 608 144
rect 651 141 653 144
rect 969 128 971 135
rect 993 128 995 135
rect 1025 134 1027 137
rect 524 109 526 116
rect 519 105 526 109
rect 520 94 522 105
rect 532 97 534 116
rect 562 108 564 116
rect 606 108 608 116
rect 556 106 564 108
rect 600 106 608 108
rect 556 94 558 106
rect 564 94 566 103
rect 600 94 602 106
rect 608 94 610 103
rect 651 94 653 116
rect 1078 130 1080 145
rect 1025 96 1027 114
rect 969 84 971 88
rect 993 84 995 88
rect 520 81 522 84
rect 556 81 558 84
rect 564 81 566 84
rect 600 81 602 84
rect 608 81 610 84
rect 651 81 653 84
rect 1025 83 1027 86
<< polycontact >>
rect 813 1086 817 1090
rect 953 1086 957 1090
rect 813 1031 817 1035
rect 882 1060 886 1064
rect 1088 1086 1092 1090
rect 893 1049 897 1053
rect 953 1031 957 1035
rect 1022 1060 1026 1064
rect 1226 1085 1230 1089
rect 1033 1049 1037 1053
rect 1088 1031 1092 1035
rect 1157 1060 1161 1064
rect 1168 1049 1172 1053
rect 1226 1030 1230 1034
rect 1295 1059 1299 1063
rect 1306 1048 1310 1052
rect 485 978 489 982
rect 498 970 502 974
rect 509 978 513 982
rect 521 970 526 975
rect 536 970 540 974
rect 565 970 570 975
rect 617 975 621 980
rect 580 970 584 974
rect 740 959 744 963
rect 750 952 754 956
rect 782 958 786 962
rect 1175 959 1179 963
rect 1004 937 1008 941
rect 1175 904 1179 908
rect 1244 933 1248 937
rect 1255 922 1259 926
rect 489 880 493 884
rect 502 872 506 876
rect 513 880 517 884
rect 525 872 530 877
rect 540 872 544 876
rect 569 872 574 877
rect 621 877 625 882
rect 584 872 588 876
rect 740 885 744 889
rect 750 878 754 882
rect 782 884 786 888
rect 913 897 917 901
rect 926 897 930 901
rect 946 897 950 901
rect 973 897 977 901
rect 996 897 1000 901
rect 1370 884 1374 888
rect 1383 876 1387 880
rect 1394 884 1398 888
rect 1406 876 1411 881
rect 1421 876 1425 880
rect 1450 876 1455 881
rect 1502 881 1506 886
rect 1465 876 1469 880
rect 1582 885 1586 889
rect 1034 846 1038 850
rect 740 816 744 820
rect 750 809 754 813
rect 782 815 786 819
rect 899 819 903 823
rect 923 819 927 823
rect 944 819 948 823
rect 961 819 965 823
rect 979 820 983 824
rect 494 782 498 786
rect 507 774 511 778
rect 518 782 522 786
rect 530 774 535 779
rect 545 774 549 778
rect 574 774 579 779
rect 626 779 630 784
rect 589 774 593 778
rect 1071 818 1075 822
rect 1018 788 1022 792
rect 1368 784 1372 788
rect 1381 776 1385 780
rect 1392 784 1396 788
rect 1404 776 1409 781
rect 1419 776 1423 780
rect 1448 776 1453 781
rect 1500 781 1504 786
rect 1463 776 1467 780
rect 1586 782 1590 786
rect 740 742 744 746
rect 750 735 754 739
rect 782 741 786 745
rect 1173 726 1177 730
rect 1000 699 1004 703
rect 501 682 505 686
rect 514 674 518 678
rect 525 682 529 686
rect 537 674 542 679
rect 552 674 556 678
rect 581 674 586 679
rect 633 679 637 684
rect 596 674 600 678
rect 1173 671 1177 675
rect 1242 700 1246 704
rect 1253 689 1257 693
rect 1367 677 1371 681
rect 926 659 930 663
rect 939 659 943 663
rect 959 659 963 663
rect 986 659 990 663
rect 1380 669 1384 673
rect 1391 677 1395 681
rect 1403 669 1408 674
rect 1418 669 1422 673
rect 1447 669 1452 674
rect 1499 674 1503 679
rect 1462 669 1466 673
rect 1588 683 1592 687
rect 1030 608 1034 612
rect 1176 602 1180 606
rect 912 581 916 585
rect 512 568 516 572
rect 525 560 529 564
rect 536 568 540 572
rect 548 560 553 565
rect 563 560 567 564
rect 592 560 597 565
rect 644 565 648 570
rect 607 560 611 564
rect 936 581 940 585
rect 957 581 961 585
rect 974 581 978 585
rect 1067 580 1071 584
rect 1014 550 1018 554
rect 1176 547 1180 551
rect 1245 576 1249 580
rect 1367 573 1371 577
rect 1256 565 1260 569
rect 1380 565 1384 569
rect 1391 573 1395 577
rect 1403 565 1408 570
rect 1418 565 1422 569
rect 1447 565 1452 570
rect 1499 570 1503 575
rect 1462 565 1466 569
rect 1584 581 1588 585
rect 1005 472 1009 476
rect 504 459 508 463
rect 517 451 521 455
rect 528 459 532 463
rect 540 451 545 456
rect 555 451 559 455
rect 584 451 589 456
rect 636 456 640 461
rect 599 451 603 455
rect 1170 454 1174 458
rect 958 432 962 436
rect 971 432 975 436
rect 991 432 995 436
rect 1367 458 1371 462
rect 1380 450 1384 454
rect 1391 458 1395 462
rect 1403 450 1408 455
rect 1418 450 1422 454
rect 1447 450 1452 455
rect 1499 455 1503 460
rect 1462 450 1466 454
rect 1581 462 1585 466
rect 1170 399 1174 403
rect 1239 428 1243 432
rect 1250 417 1254 421
rect 1035 381 1039 385
rect 944 354 948 358
rect 968 354 972 358
rect 989 354 993 358
rect 509 334 513 338
rect 522 326 526 330
rect 533 334 537 338
rect 545 326 550 331
rect 560 326 564 330
rect 589 326 594 331
rect 641 331 645 336
rect 604 326 608 330
rect 1072 353 1076 357
rect 1019 323 1023 327
rect 1007 249 1011 253
rect 525 223 529 227
rect 538 215 542 219
rect 549 223 553 227
rect 561 215 566 220
rect 576 215 580 219
rect 605 215 610 220
rect 657 220 661 225
rect 620 215 624 219
rect 979 209 983 213
rect 992 209 996 213
rect 1037 158 1041 162
rect 965 131 969 135
rect 989 131 993 135
rect 515 105 519 109
rect 528 97 532 101
rect 539 105 543 109
rect 551 97 556 102
rect 566 97 570 101
rect 595 97 600 102
rect 647 102 651 107
rect 610 97 614 101
rect 1074 130 1078 134
rect 1021 100 1025 104
<< metal1 >>
rect 811 1115 839 1118
rect 951 1115 979 1118
rect 1086 1115 1114 1118
rect 812 1109 815 1115
rect 836 1114 839 1115
rect 836 1111 907 1114
rect 795 1085 798 1088
rect 803 1086 813 1089
rect 821 1089 824 1097
rect 851 1105 854 1111
rect 870 1105 873 1111
rect 952 1109 955 1115
rect 976 1114 979 1115
rect 976 1111 1047 1114
rect 821 1086 842 1089
rect 821 1083 824 1086
rect 812 1073 815 1077
rect 806 1071 830 1073
rect 806 1070 824 1071
rect 829 1070 830 1071
rect 839 1063 842 1086
rect 880 1105 900 1108
rect 880 1099 883 1105
rect 897 1099 900 1105
rect 861 1078 864 1081
rect 861 1075 879 1078
rect 935 1085 938 1088
rect 943 1086 953 1089
rect 961 1089 964 1097
rect 991 1105 994 1111
rect 1010 1105 1013 1111
rect 1087 1109 1090 1115
rect 1111 1114 1114 1115
rect 1224 1114 1252 1117
rect 1111 1111 1182 1114
rect 961 1086 982 1089
rect 961 1083 964 1086
rect 889 1068 892 1075
rect 952 1073 955 1077
rect 946 1071 970 1073
rect 946 1070 964 1071
rect 889 1065 906 1068
rect 811 1062 830 1063
rect 806 1060 830 1062
rect 839 1060 882 1063
rect 812 1054 815 1060
rect 903 1054 906 1065
rect 969 1070 970 1071
rect 979 1063 982 1086
rect 1020 1105 1040 1108
rect 1020 1099 1023 1105
rect 1037 1099 1040 1105
rect 1001 1078 1004 1081
rect 1001 1075 1019 1078
rect 1070 1085 1073 1088
rect 1078 1086 1088 1089
rect 1096 1089 1099 1097
rect 1126 1105 1129 1111
rect 1145 1105 1148 1111
rect 1225 1108 1228 1114
rect 1249 1113 1252 1114
rect 1249 1110 1320 1113
rect 1096 1086 1117 1089
rect 1096 1083 1099 1086
rect 1029 1068 1032 1075
rect 1087 1073 1090 1077
rect 1081 1071 1105 1073
rect 1081 1070 1099 1071
rect 1029 1065 1046 1068
rect 951 1062 970 1063
rect 946 1060 970 1062
rect 979 1060 1022 1063
rect 952 1054 955 1060
rect 1043 1054 1046 1065
rect 1104 1070 1105 1071
rect 1114 1063 1117 1086
rect 1155 1105 1175 1108
rect 1155 1099 1158 1105
rect 1172 1099 1175 1105
rect 1136 1078 1139 1081
rect 1136 1075 1154 1078
rect 1208 1084 1211 1087
rect 1216 1085 1226 1088
rect 1234 1088 1237 1096
rect 1264 1104 1267 1110
rect 1283 1104 1286 1110
rect 1234 1085 1255 1088
rect 1234 1082 1237 1085
rect 1164 1068 1167 1075
rect 1225 1072 1228 1076
rect 1219 1070 1243 1072
rect 1219 1069 1237 1070
rect 1164 1065 1181 1068
rect 1086 1062 1105 1063
rect 1081 1060 1105 1062
rect 1114 1060 1157 1063
rect 1087 1054 1090 1060
rect 1178 1054 1181 1065
rect 1242 1069 1243 1070
rect 1252 1062 1255 1085
rect 1293 1104 1313 1107
rect 1293 1098 1296 1104
rect 1310 1098 1313 1104
rect 1274 1077 1277 1080
rect 1274 1074 1292 1077
rect 1302 1067 1305 1074
rect 1302 1064 1319 1067
rect 1224 1061 1243 1062
rect 1219 1059 1243 1061
rect 1252 1059 1295 1062
rect 868 1049 893 1052
rect 903 1050 916 1054
rect 868 1047 871 1049
rect 795 1031 798 1034
rect 803 1031 813 1034
rect 821 1034 824 1042
rect 833 1044 871 1047
rect 903 1046 906 1050
rect 833 1034 836 1044
rect 874 1043 906 1046
rect 874 1040 877 1043
rect 821 1031 836 1034
rect 821 1028 824 1031
rect 483 1020 636 1024
rect 873 1037 879 1040
rect 489 1014 493 1020
rect 527 1014 531 1020
rect 571 1014 575 1020
rect 616 1014 620 1020
rect 812 1018 815 1022
rect 833 1021 838 1024
rect 851 1024 854 1028
rect 898 1024 901 1028
rect 843 1021 907 1024
rect 833 1018 836 1021
rect 806 1015 836 1018
rect 539 989 552 1014
rect 583 989 596 1014
rect 912 1010 916 1050
rect 1008 1049 1033 1052
rect 1043 1050 1055 1054
rect 1008 1047 1011 1049
rect 935 1031 938 1034
rect 943 1031 953 1034
rect 961 1034 964 1042
rect 973 1044 1011 1047
rect 1043 1046 1046 1050
rect 973 1034 976 1044
rect 1014 1043 1046 1046
rect 1014 1040 1017 1043
rect 961 1031 976 1034
rect 961 1028 964 1031
rect 1013 1037 1019 1040
rect 952 1018 955 1022
rect 973 1021 978 1024
rect 991 1024 994 1028
rect 1038 1024 1041 1028
rect 983 1021 1047 1024
rect 973 1018 976 1021
rect 946 1015 976 1018
rect 1051 1009 1055 1050
rect 1143 1049 1168 1052
rect 1178 1050 1189 1054
rect 1143 1047 1146 1049
rect 1070 1031 1073 1034
rect 1078 1031 1088 1034
rect 1096 1034 1099 1042
rect 1108 1044 1146 1047
rect 1178 1046 1181 1050
rect 1108 1034 1111 1044
rect 1149 1043 1181 1046
rect 1149 1040 1152 1043
rect 1096 1031 1111 1034
rect 1096 1028 1099 1031
rect 1148 1037 1154 1040
rect 1087 1018 1090 1022
rect 1108 1021 1113 1024
rect 1126 1024 1129 1028
rect 1173 1024 1176 1028
rect 1118 1021 1182 1024
rect 1108 1018 1111 1021
rect 1081 1015 1111 1018
rect 1185 1010 1189 1050
rect 1225 1053 1228 1059
rect 1316 1053 1319 1064
rect 1281 1048 1306 1051
rect 1316 1049 1331 1053
rect 1281 1046 1284 1048
rect 1208 1030 1211 1033
rect 1216 1030 1226 1033
rect 1234 1033 1237 1041
rect 1246 1043 1284 1046
rect 1316 1045 1319 1049
rect 1246 1033 1249 1043
rect 1287 1042 1319 1045
rect 1287 1039 1290 1042
rect 1234 1030 1249 1033
rect 1234 1027 1237 1030
rect 1286 1036 1292 1039
rect 1225 1017 1228 1021
rect 1246 1020 1251 1023
rect 1264 1023 1267 1027
rect 1311 1023 1314 1027
rect 1256 1020 1320 1023
rect 1246 1017 1249 1020
rect 1219 1014 1249 1017
rect 1327 1011 1331 1049
rect 1051 1005 1058 1009
rect 1182 1006 1189 1010
rect 731 990 802 993
rect 478 978 485 982
rect 489 970 498 974
rect 505 967 509 989
rect 513 978 514 982
rect 549 980 552 989
rect 593 980 596 989
rect 549 975 561 980
rect 593 975 617 980
rect 624 979 628 989
rect 739 984 743 990
rect 757 984 761 990
rect 513 973 521 975
rect 518 970 521 973
rect 540 970 541 974
rect 549 967 552 975
rect 557 970 565 975
rect 584 970 585 974
rect 593 967 596 975
rect 624 974 637 979
rect 624 967 628 974
rect 781 984 784 990
rect 1173 988 1201 991
rect 1174 982 1177 988
rect 1198 987 1201 988
rect 1198 984 1269 987
rect 996 977 1024 980
rect 497 957 509 967
rect 541 957 552 967
rect 585 957 596 967
rect 748 969 751 972
rect 748 966 761 969
rect 731 959 740 963
rect 758 962 761 966
rect 790 962 793 972
rect 1003 971 1006 977
rect 758 958 782 962
rect 790 959 802 962
rect 485 952 489 957
rect 521 952 525 957
rect 565 952 569 957
rect 616 952 620 957
rect 731 952 750 956
rect 484 948 628 952
rect 758 949 761 958
rect 790 954 793 959
rect 1157 958 1160 961
rect 1165 959 1175 962
rect 1183 962 1186 970
rect 1213 978 1216 984
rect 1232 978 1235 984
rect 1183 959 1204 962
rect 1183 956 1186 959
rect 739 930 742 936
rect 781 930 784 947
rect 1012 941 1015 951
rect 1174 946 1177 950
rect 1168 944 1192 946
rect 1168 943 1186 944
rect 996 937 1004 941
rect 1012 938 1024 941
rect 1012 933 1015 938
rect 1191 943 1192 944
rect 1201 936 1204 959
rect 1242 978 1262 981
rect 1242 972 1245 978
rect 1259 972 1262 978
rect 1223 951 1226 954
rect 1223 948 1241 951
rect 1251 941 1254 948
rect 1251 938 1268 941
rect 1173 935 1192 936
rect 1168 933 1192 935
rect 1201 933 1244 936
rect 731 927 784 930
rect 487 922 640 926
rect 1174 927 1177 933
rect 1265 927 1268 938
rect 493 916 497 922
rect 531 916 535 922
rect 575 916 579 922
rect 620 916 624 922
rect 731 916 802 919
rect 543 891 556 916
rect 587 891 600 916
rect 739 910 743 916
rect 757 910 761 916
rect 781 910 784 916
rect 1003 915 1006 923
rect 1230 922 1255 925
rect 1265 923 1278 927
rect 1368 926 1521 930
rect 1230 920 1233 922
rect 996 912 1006 915
rect 1018 909 1021 911
rect 748 895 751 898
rect 748 892 761 895
rect 482 880 489 884
rect 493 872 502 876
rect 509 869 513 891
rect 517 880 518 884
rect 553 882 556 891
rect 597 882 600 891
rect 553 877 565 882
rect 597 877 621 882
rect 628 881 632 891
rect 731 885 740 889
rect 758 888 761 892
rect 790 888 793 898
rect 910 897 913 901
rect 930 897 936 901
rect 943 897 946 901
rect 970 897 973 901
rect 993 897 996 901
rect 1003 900 1007 901
rect 1003 896 1014 900
rect 1003 894 1007 896
rect 758 884 782 888
rect 790 885 802 888
rect 517 875 525 877
rect 522 872 525 875
rect 544 872 545 876
rect 553 869 556 877
rect 561 872 569 877
rect 588 872 589 876
rect 597 869 600 877
rect 628 876 641 881
rect 731 878 750 882
rect 628 869 632 876
rect 758 875 761 884
rect 790 880 793 885
rect 501 859 513 869
rect 545 859 556 869
rect 589 859 600 869
rect 489 854 493 859
rect 525 854 529 859
rect 569 854 573 859
rect 620 854 624 859
rect 739 856 742 862
rect 781 856 784 873
rect 488 850 632 854
rect 731 853 784 856
rect 731 847 802 850
rect 739 841 743 847
rect 757 841 761 847
rect 781 841 784 847
rect 912 844 916 853
rect 927 852 932 853
rect 945 852 949 854
rect 927 847 949 852
rect 953 852 957 854
rect 972 852 976 854
rect 953 847 976 852
rect 980 852 984 854
rect 995 852 999 854
rect 980 847 999 852
rect 907 840 925 844
rect 492 824 645 828
rect 748 826 751 829
rect 498 818 502 824
rect 536 818 540 824
rect 580 818 584 824
rect 625 818 629 824
rect 748 823 761 826
rect 548 793 561 818
rect 592 793 605 818
rect 731 816 740 820
rect 758 819 761 823
rect 790 819 793 829
rect 896 819 899 823
rect 758 815 782 819
rect 790 816 802 819
rect 906 816 910 825
rect 731 809 750 813
rect 758 806 761 815
rect 790 811 793 816
rect 487 782 494 786
rect 498 774 507 778
rect 514 771 518 793
rect 522 782 523 786
rect 558 784 561 793
rect 602 784 605 793
rect 558 779 570 784
rect 602 779 626 784
rect 633 783 637 793
rect 739 787 742 793
rect 781 787 784 804
rect 731 784 784 787
rect 522 777 530 779
rect 527 774 530 777
rect 549 774 550 778
rect 558 771 561 779
rect 566 774 574 779
rect 593 774 594 778
rect 602 771 605 779
rect 633 778 646 783
rect 633 771 637 778
rect 731 773 802 776
rect 506 761 518 771
rect 550 761 561 771
rect 594 761 605 771
rect 739 767 743 773
rect 757 767 761 773
rect 494 756 498 761
rect 530 756 534 761
rect 574 756 578 761
rect 625 756 629 761
rect 493 752 637 756
rect 781 767 784 773
rect 898 771 902 776
rect 913 771 917 840
rect 920 819 923 823
rect 930 816 934 847
rect 958 840 962 847
rect 985 840 989 847
rect 1010 845 1014 896
rect 1017 850 1021 909
rect 1026 907 1054 910
rect 1033 901 1036 907
rect 1157 904 1160 907
rect 1165 904 1175 907
rect 1183 907 1186 915
rect 1195 917 1233 920
rect 1265 919 1268 923
rect 1195 907 1198 917
rect 1236 916 1268 919
rect 1236 913 1239 916
rect 1183 904 1198 907
rect 1183 901 1186 904
rect 1235 910 1241 913
rect 1174 891 1177 895
rect 1195 894 1200 897
rect 1213 897 1216 901
rect 1260 897 1263 901
rect 1205 894 1269 897
rect 1195 891 1198 894
rect 1168 888 1198 891
rect 1274 883 1278 923
rect 1374 920 1378 926
rect 1412 920 1416 926
rect 1456 920 1460 926
rect 1501 920 1505 926
rect 1574 925 1602 928
rect 1424 895 1437 920
rect 1468 895 1481 920
rect 1581 919 1584 925
rect 1363 884 1370 888
rect 1374 876 1383 880
rect 1390 873 1394 895
rect 1398 884 1399 888
rect 1434 886 1437 895
rect 1478 886 1481 895
rect 1434 881 1446 886
rect 1478 881 1502 886
rect 1509 885 1513 895
rect 1590 889 1593 899
rect 1574 885 1582 889
rect 1590 886 1602 889
rect 1398 879 1406 881
rect 1403 876 1406 879
rect 1425 876 1426 880
rect 1434 873 1437 881
rect 1442 876 1450 881
rect 1469 876 1470 880
rect 1478 873 1481 881
rect 1509 880 1522 885
rect 1590 881 1593 886
rect 1509 873 1513 880
rect 1017 846 1034 850
rect 1042 849 1045 861
rect 1382 863 1394 873
rect 1426 863 1437 873
rect 1470 863 1481 873
rect 1581 863 1584 871
rect 1057 856 1098 859
rect 1370 858 1374 863
rect 1406 858 1410 863
rect 1450 858 1454 863
rect 1501 858 1505 863
rect 1574 860 1584 863
rect 1057 849 1060 856
rect 1063 849 1091 852
rect 1042 846 1060 849
rect 951 836 962 840
rect 968 836 989 840
rect 1002 843 1014 845
rect 1046 843 1050 846
rect 1002 841 1050 843
rect 941 819 944 823
rect 951 816 955 836
rect 958 819 961 823
rect 968 816 972 836
rect 1002 824 1006 841
rect 1010 839 1050 841
rect 1070 843 1073 849
rect 1010 828 1038 831
rect 976 820 979 824
rect 986 820 1006 824
rect 986 817 990 820
rect 1002 792 1006 820
rect 1017 822 1020 828
rect 1026 792 1029 802
rect 1041 819 1071 822
rect 1041 792 1044 819
rect 1063 818 1071 819
rect 1079 821 1082 833
rect 1095 821 1098 856
rect 1369 854 1513 858
rect 1366 826 1519 830
rect 1079 818 1098 821
rect 1372 820 1376 826
rect 1410 820 1414 826
rect 1454 820 1458 826
rect 1499 820 1503 826
rect 1578 822 1606 825
rect 1422 795 1435 820
rect 1466 795 1479 820
rect 1585 816 1588 822
rect 1002 788 1018 792
rect 1026 789 1044 792
rect 1026 784 1029 789
rect 1361 784 1368 788
rect 922 771 926 776
rect 943 771 947 776
rect 960 771 964 776
rect 978 771 982 777
rect 898 768 982 771
rect 1372 776 1381 780
rect 1017 766 1020 774
rect 1388 773 1392 795
rect 1396 784 1397 788
rect 1432 786 1435 795
rect 1476 786 1479 795
rect 1432 781 1444 786
rect 1476 781 1500 786
rect 1507 785 1511 795
rect 1594 786 1597 796
rect 1396 779 1404 781
rect 1401 776 1404 779
rect 1423 776 1424 780
rect 1432 773 1435 781
rect 1440 776 1448 781
rect 1467 776 1468 780
rect 1476 773 1479 781
rect 1507 780 1520 785
rect 1578 782 1586 786
rect 1594 783 1606 786
rect 1507 773 1511 780
rect 1594 778 1597 783
rect 1006 763 1020 766
rect 1380 763 1392 773
rect 1424 763 1435 773
rect 1468 763 1479 773
rect 1368 758 1372 763
rect 1404 758 1408 763
rect 1448 758 1452 763
rect 1499 758 1503 763
rect 1585 760 1588 768
rect 1171 755 1199 758
rect 748 752 751 755
rect 748 749 761 752
rect 731 742 740 746
rect 758 745 761 749
rect 790 745 793 755
rect 1172 749 1175 755
rect 1196 754 1199 755
rect 1367 754 1511 758
rect 1578 757 1588 760
rect 1196 751 1267 754
rect 758 741 782 745
rect 790 742 802 745
rect 731 735 750 739
rect 758 732 761 741
rect 790 737 793 742
rect 992 739 1020 742
rect 499 724 652 728
rect 505 718 509 724
rect 543 718 547 724
rect 587 718 591 724
rect 632 718 636 724
rect 999 733 1002 739
rect 555 693 568 718
rect 599 693 612 718
rect 739 713 742 719
rect 781 713 784 730
rect 1155 725 1158 728
rect 1163 726 1173 729
rect 1181 729 1184 737
rect 1211 745 1214 751
rect 1230 745 1233 751
rect 1181 726 1202 729
rect 1181 723 1184 726
rect 1172 713 1175 717
rect 731 710 784 713
rect 1008 703 1011 713
rect 1166 711 1190 713
rect 1166 710 1184 711
rect 992 699 1000 703
rect 1008 700 1020 703
rect 1189 710 1190 711
rect 1199 703 1202 726
rect 1240 745 1260 748
rect 1240 739 1243 745
rect 1257 739 1260 745
rect 1221 718 1224 721
rect 1221 715 1239 718
rect 1580 723 1608 726
rect 1365 719 1518 723
rect 1249 708 1252 715
rect 1371 713 1375 719
rect 1409 713 1413 719
rect 1453 713 1457 719
rect 1498 713 1502 719
rect 1587 717 1590 723
rect 1249 705 1266 708
rect 1171 702 1190 703
rect 1166 700 1190 702
rect 1199 700 1242 703
rect 1008 695 1011 700
rect 494 682 501 686
rect 505 674 514 678
rect 521 671 525 693
rect 529 682 530 686
rect 565 684 568 693
rect 609 684 612 693
rect 565 679 577 684
rect 609 679 633 684
rect 640 683 644 693
rect 1172 694 1175 700
rect 1263 694 1266 705
rect 529 677 537 679
rect 534 674 537 677
rect 556 674 557 678
rect 565 671 568 679
rect 573 674 581 679
rect 600 674 601 678
rect 609 671 612 679
rect 640 678 653 683
rect 640 671 644 678
rect 999 677 1002 685
rect 1228 689 1253 692
rect 1263 690 1276 694
rect 1228 687 1231 689
rect 992 674 1002 677
rect 1014 671 1017 673
rect 513 661 525 671
rect 557 661 568 671
rect 601 661 612 671
rect 501 656 505 661
rect 537 656 541 661
rect 581 656 585 661
rect 632 656 636 661
rect 923 659 926 663
rect 943 659 949 663
rect 956 659 959 663
rect 983 659 986 663
rect 500 652 644 656
rect 510 610 663 614
rect 516 604 520 610
rect 554 604 558 610
rect 598 604 602 610
rect 643 604 647 610
rect 925 606 929 615
rect 940 614 945 615
rect 958 614 962 616
rect 940 609 962 614
rect 966 614 970 616
rect 985 614 989 616
rect 966 609 989 614
rect 993 614 997 616
rect 993 609 1002 614
rect 566 579 579 604
rect 610 579 623 604
rect 920 602 938 606
rect 909 581 912 585
rect 505 568 512 572
rect 516 560 525 564
rect 532 557 536 579
rect 540 568 541 572
rect 576 570 579 579
rect 620 570 623 579
rect 576 565 588 570
rect 620 565 644 570
rect 651 569 655 579
rect 919 578 923 587
rect 540 563 548 565
rect 545 560 548 563
rect 567 560 568 564
rect 576 557 579 565
rect 584 560 592 565
rect 611 560 612 564
rect 620 557 623 565
rect 651 564 664 569
rect 651 557 655 564
rect 524 547 536 557
rect 568 547 579 557
rect 612 547 623 557
rect 512 542 516 547
rect 548 542 552 547
rect 592 542 596 547
rect 643 542 647 547
rect 511 538 655 542
rect 911 533 915 538
rect 926 533 930 602
rect 933 581 936 585
rect 943 578 947 609
rect 971 602 975 609
rect 998 605 1002 609
rect 1013 612 1017 671
rect 1022 669 1050 672
rect 1155 671 1158 674
rect 1163 671 1173 674
rect 1181 674 1184 682
rect 1193 684 1231 687
rect 1263 686 1266 690
rect 1193 674 1196 684
rect 1234 683 1266 686
rect 1234 680 1237 683
rect 1181 671 1196 674
rect 1029 663 1032 669
rect 1181 668 1184 671
rect 1233 677 1239 680
rect 1172 658 1175 662
rect 1193 661 1198 664
rect 1211 664 1214 668
rect 1258 664 1261 668
rect 1203 661 1267 664
rect 1193 658 1196 661
rect 1166 655 1196 658
rect 1272 650 1276 690
rect 1421 688 1434 713
rect 1465 688 1478 713
rect 1360 677 1367 681
rect 1371 669 1380 673
rect 1387 666 1391 688
rect 1395 677 1396 681
rect 1431 679 1434 688
rect 1475 679 1478 688
rect 1431 674 1443 679
rect 1475 674 1499 679
rect 1506 678 1510 688
rect 1596 687 1599 697
rect 1580 683 1588 687
rect 1596 684 1608 687
rect 1596 679 1599 684
rect 1395 672 1403 674
rect 1400 669 1403 672
rect 1422 669 1423 673
rect 1431 666 1434 674
rect 1439 669 1447 674
rect 1466 669 1467 673
rect 1475 666 1478 674
rect 1506 673 1519 678
rect 1506 666 1510 673
rect 1379 656 1391 666
rect 1423 656 1434 666
rect 1467 656 1478 666
rect 1587 661 1590 669
rect 1580 658 1590 661
rect 1367 651 1371 656
rect 1403 651 1407 656
rect 1447 651 1451 656
rect 1498 651 1502 656
rect 1366 647 1510 651
rect 1174 631 1202 634
rect 1013 608 1030 612
rect 1038 611 1041 623
rect 1175 625 1178 631
rect 1199 630 1202 631
rect 1199 627 1270 630
rect 1053 618 1094 621
rect 1053 611 1056 618
rect 1059 611 1087 614
rect 1038 608 1056 611
rect 1042 605 1046 608
rect 964 598 975 602
rect 981 601 1046 605
rect 1066 605 1069 611
rect 954 581 957 585
rect 964 578 968 598
rect 971 581 974 585
rect 981 578 985 601
rect 998 554 1002 601
rect 1006 590 1034 593
rect 1013 584 1016 590
rect 1022 554 1025 564
rect 1037 581 1067 584
rect 1037 554 1040 581
rect 1059 580 1067 581
rect 1075 583 1078 595
rect 1091 583 1094 618
rect 1158 601 1161 604
rect 1166 602 1176 605
rect 1184 605 1187 613
rect 1214 621 1217 627
rect 1233 621 1236 627
rect 1184 602 1205 605
rect 1184 599 1187 602
rect 1175 589 1178 593
rect 1169 587 1193 589
rect 1169 586 1187 587
rect 1075 580 1094 583
rect 1192 586 1193 587
rect 1202 579 1205 602
rect 1243 621 1263 624
rect 1576 621 1604 624
rect 1243 615 1246 621
rect 1260 615 1263 621
rect 1365 615 1518 619
rect 1583 615 1586 621
rect 1224 594 1227 597
rect 1224 591 1242 594
rect 1371 609 1375 615
rect 1409 609 1413 615
rect 1453 609 1457 615
rect 1498 609 1502 615
rect 1252 584 1255 591
rect 1421 584 1434 609
rect 1465 584 1478 609
rect 1592 585 1595 595
rect 1252 581 1269 584
rect 1174 578 1193 579
rect 1169 576 1193 578
rect 1202 576 1245 579
rect 1175 570 1178 576
rect 1266 570 1269 581
rect 1360 573 1367 577
rect 1231 565 1256 568
rect 1266 566 1279 570
rect 1231 563 1234 565
rect 998 550 1014 554
rect 1022 551 1040 554
rect 1022 546 1025 551
rect 1158 547 1161 550
rect 1166 547 1176 550
rect 1184 550 1187 558
rect 1196 560 1234 563
rect 1266 562 1269 566
rect 1196 550 1199 560
rect 1237 559 1269 562
rect 1237 556 1240 559
rect 1184 547 1199 550
rect 935 533 939 538
rect 956 533 960 538
rect 973 533 977 538
rect 1184 544 1187 547
rect 1236 553 1242 556
rect 911 530 978 533
rect 1013 528 1016 536
rect 1175 534 1178 538
rect 1196 537 1201 540
rect 1214 540 1217 544
rect 1261 540 1264 544
rect 1206 537 1270 540
rect 1196 534 1199 537
rect 1169 531 1199 534
rect 1002 525 1016 528
rect 1275 526 1279 566
rect 1371 565 1380 569
rect 1387 562 1391 584
rect 1395 573 1396 577
rect 1431 575 1434 584
rect 1475 575 1478 584
rect 1431 570 1443 575
rect 1475 570 1499 575
rect 1506 574 1510 584
rect 1576 581 1584 585
rect 1592 582 1604 585
rect 1592 577 1595 582
rect 1395 568 1403 570
rect 1400 565 1403 568
rect 1422 565 1423 569
rect 1431 562 1434 570
rect 1439 565 1447 570
rect 1466 565 1467 569
rect 1475 562 1478 570
rect 1506 569 1519 574
rect 1506 562 1510 569
rect 1379 552 1391 562
rect 1423 552 1434 562
rect 1467 552 1478 562
rect 1583 559 1586 567
rect 1576 556 1586 559
rect 1367 547 1371 552
rect 1403 547 1407 552
rect 1447 547 1451 552
rect 1498 547 1502 552
rect 1366 543 1510 547
rect 997 512 1025 515
rect 1004 506 1007 512
rect 502 501 655 505
rect 508 495 512 501
rect 546 495 550 501
rect 590 495 594 501
rect 635 495 639 501
rect 558 470 571 495
rect 602 470 615 495
rect 1365 500 1518 504
rect 1573 502 1601 505
rect 1371 494 1375 500
rect 1409 494 1413 500
rect 1453 494 1457 500
rect 1498 494 1502 500
rect 1580 496 1583 502
rect 1013 476 1016 486
rect 1168 483 1196 486
rect 1169 477 1172 483
rect 1193 482 1196 483
rect 1193 479 1264 482
rect 997 472 1005 476
rect 1013 473 1025 476
rect 497 459 504 463
rect 508 451 517 455
rect 524 448 528 470
rect 532 459 533 463
rect 568 461 571 470
rect 612 461 615 470
rect 568 456 580 461
rect 612 456 636 461
rect 643 460 647 470
rect 1013 468 1016 473
rect 532 454 540 456
rect 537 451 540 454
rect 559 451 560 455
rect 568 448 571 456
rect 576 451 584 456
rect 603 451 604 455
rect 612 448 615 456
rect 643 455 656 460
rect 643 448 647 455
rect 1004 450 1007 458
rect 1152 453 1155 456
rect 1160 454 1170 457
rect 1178 457 1181 465
rect 1208 473 1211 479
rect 1227 473 1230 479
rect 1178 454 1199 457
rect 1178 451 1181 454
rect 516 438 528 448
rect 560 438 571 448
rect 604 438 615 448
rect 997 447 1007 450
rect 1019 444 1022 446
rect 504 433 508 438
rect 540 433 544 438
rect 584 433 588 438
rect 635 433 639 438
rect 503 429 647 433
rect 955 432 958 436
rect 975 432 981 436
rect 988 432 991 436
rect 507 376 660 380
rect 957 379 961 388
rect 972 387 977 388
rect 990 387 994 389
rect 972 382 994 387
rect 998 387 1002 389
rect 998 385 1004 387
rect 1018 385 1022 444
rect 1027 442 1055 445
rect 1034 436 1037 442
rect 1169 441 1172 445
rect 1163 439 1187 441
rect 1163 438 1181 439
rect 1186 438 1187 439
rect 1196 431 1199 454
rect 1237 473 1257 476
rect 1237 467 1240 473
rect 1254 467 1257 473
rect 1421 469 1434 494
rect 1465 469 1478 494
rect 1218 446 1221 449
rect 1218 443 1236 446
rect 1360 458 1367 462
rect 1371 450 1380 454
rect 1387 447 1391 469
rect 1395 458 1396 462
rect 1431 460 1434 469
rect 1475 460 1478 469
rect 1431 455 1443 460
rect 1475 455 1499 460
rect 1506 459 1510 469
rect 1589 466 1592 476
rect 1573 462 1581 466
rect 1589 463 1601 466
rect 1395 453 1403 455
rect 1400 450 1403 453
rect 1422 450 1423 454
rect 1431 447 1434 455
rect 1439 450 1447 455
rect 1466 450 1467 454
rect 1475 447 1478 455
rect 1506 454 1519 459
rect 1589 458 1592 463
rect 1506 447 1510 454
rect 1246 436 1249 443
rect 1379 437 1391 447
rect 1423 437 1434 447
rect 1467 437 1478 447
rect 1580 440 1583 448
rect 1573 437 1583 440
rect 1246 433 1263 436
rect 1168 430 1187 431
rect 1163 428 1187 430
rect 1196 428 1239 431
rect 1169 422 1172 428
rect 1260 422 1263 433
rect 1367 432 1371 437
rect 1403 432 1407 437
rect 1447 432 1451 437
rect 1498 432 1502 437
rect 1366 428 1510 432
rect 1225 417 1250 420
rect 1260 418 1273 422
rect 1225 415 1228 417
rect 1152 399 1155 402
rect 1160 399 1170 402
rect 1178 402 1181 410
rect 1190 412 1228 415
rect 1260 414 1263 418
rect 1190 402 1193 412
rect 1231 411 1263 414
rect 1231 408 1234 411
rect 1178 399 1193 402
rect 1178 396 1181 399
rect 998 382 1006 385
rect 513 370 517 376
rect 551 370 555 376
rect 595 370 599 376
rect 640 370 644 376
rect 952 375 970 379
rect 563 345 576 370
rect 607 345 620 370
rect 941 354 944 358
rect 951 351 955 360
rect 502 334 509 338
rect 513 326 522 330
rect 529 323 533 345
rect 537 334 538 338
rect 573 336 576 345
rect 617 336 620 345
rect 573 331 585 336
rect 617 331 641 336
rect 648 335 652 345
rect 537 329 545 331
rect 542 326 545 329
rect 564 326 565 330
rect 573 323 576 331
rect 581 326 589 331
rect 608 326 609 330
rect 617 323 620 331
rect 648 330 661 335
rect 648 323 652 330
rect 521 313 533 323
rect 565 313 576 323
rect 609 313 620 323
rect 509 308 513 313
rect 545 308 549 313
rect 589 308 593 313
rect 640 308 644 313
rect 508 304 652 308
rect 943 306 947 311
rect 958 306 962 375
rect 965 354 968 358
rect 975 351 979 382
rect 1002 378 1006 382
rect 1018 381 1035 385
rect 1043 384 1046 396
rect 1058 391 1099 394
rect 1058 384 1061 391
rect 1064 384 1092 387
rect 1043 381 1061 384
rect 1047 378 1051 381
rect 1002 375 1051 378
rect 996 374 1051 375
rect 1071 378 1074 384
rect 996 371 1009 374
rect 986 354 989 358
rect 996 351 1000 371
rect 1003 327 1007 371
rect 1011 363 1039 366
rect 1018 357 1021 363
rect 1027 327 1030 337
rect 1042 354 1072 357
rect 1042 327 1045 354
rect 1064 353 1072 354
rect 1080 356 1083 368
rect 1096 356 1099 391
rect 1230 405 1236 408
rect 1169 386 1172 390
rect 1190 389 1195 392
rect 1208 392 1211 396
rect 1255 392 1258 396
rect 1200 389 1264 392
rect 1190 386 1193 389
rect 1163 383 1193 386
rect 1269 378 1273 418
rect 1080 353 1099 356
rect 1003 323 1019 327
rect 1027 324 1045 327
rect 1027 319 1030 324
rect 967 306 971 311
rect 988 306 992 311
rect 943 303 1002 306
rect 1018 301 1021 309
rect 1007 298 1021 301
rect 999 289 1027 292
rect 1006 283 1009 289
rect 523 265 676 269
rect 529 259 533 265
rect 567 259 571 265
rect 611 259 615 265
rect 656 259 660 265
rect 579 234 592 259
rect 623 234 636 259
rect 1015 253 1018 263
rect 999 249 1007 253
rect 1015 250 1027 253
rect 1015 245 1018 250
rect 518 223 525 227
rect 529 215 538 219
rect 545 212 549 234
rect 553 223 554 227
rect 589 225 592 234
rect 633 225 636 234
rect 589 220 601 225
rect 633 220 657 225
rect 664 224 668 234
rect 1006 227 1009 235
rect 999 224 1009 227
rect 553 218 561 220
rect 558 215 561 218
rect 580 215 581 219
rect 589 212 592 220
rect 597 215 605 220
rect 624 215 625 219
rect 633 212 636 220
rect 664 219 677 224
rect 1021 221 1024 223
rect 664 212 668 219
rect 537 202 549 212
rect 581 202 592 212
rect 625 202 636 212
rect 976 209 979 213
rect 996 209 1002 213
rect 525 197 529 202
rect 561 197 565 202
rect 605 197 609 202
rect 656 197 660 202
rect 524 193 668 197
rect 978 156 982 165
rect 993 164 998 165
rect 993 159 999 164
rect 1020 162 1024 221
rect 1029 219 1057 222
rect 1036 213 1039 219
rect 973 152 991 156
rect 996 155 1000 159
rect 1020 158 1037 162
rect 1045 161 1048 173
rect 1060 168 1101 171
rect 1060 161 1063 168
rect 1066 161 1094 164
rect 1045 158 1063 161
rect 1049 155 1053 158
rect 513 147 666 151
rect 519 141 523 147
rect 557 141 561 147
rect 601 141 605 147
rect 646 141 650 147
rect 569 116 582 141
rect 613 116 626 141
rect 962 131 965 135
rect 972 128 976 137
rect 508 105 515 109
rect 519 97 528 101
rect 535 94 539 116
rect 543 105 544 109
rect 579 107 582 116
rect 623 107 626 116
rect 579 102 591 107
rect 623 102 647 107
rect 654 106 658 116
rect 543 100 551 102
rect 548 97 551 100
rect 570 97 571 101
rect 579 94 582 102
rect 587 97 595 102
rect 614 97 615 101
rect 623 94 626 102
rect 654 101 667 106
rect 654 94 658 101
rect 527 84 539 94
rect 571 84 582 94
rect 615 84 626 94
rect 515 79 519 84
rect 551 79 555 84
rect 595 79 599 84
rect 646 79 650 84
rect 964 83 968 88
rect 979 83 983 152
rect 996 151 1053 155
rect 1073 155 1076 161
rect 986 131 989 135
rect 996 128 1000 151
rect 1005 104 1009 151
rect 1013 140 1041 143
rect 1020 134 1023 140
rect 1029 104 1032 114
rect 1044 131 1074 134
rect 1044 104 1047 131
rect 1066 130 1074 131
rect 1082 133 1085 145
rect 1098 133 1101 168
rect 1082 130 1101 133
rect 1005 100 1021 104
rect 1029 101 1047 104
rect 1029 96 1032 101
rect 988 83 992 88
rect 964 80 1006 83
rect 514 75 658 79
rect 1020 78 1023 86
rect 1009 75 1023 78
<< m2contact >>
rect 798 1084 803 1089
rect 938 1084 943 1089
rect 1073 1084 1078 1089
rect 1211 1083 1216 1088
rect 798 1030 803 1035
rect 938 1030 943 1035
rect 1073 1030 1078 1035
rect 1211 1029 1216 1034
rect 484 970 489 975
rect 514 978 519 983
rect 513 968 518 973
rect 541 970 546 975
rect 585 970 590 975
rect 1160 957 1165 962
rect 488 872 493 877
rect 518 880 523 885
rect 517 870 522 875
rect 545 872 550 877
rect 589 872 594 877
rect 493 774 498 779
rect 523 782 528 787
rect 522 772 527 777
rect 550 774 555 779
rect 594 774 599 779
rect 1160 903 1165 908
rect 1369 876 1374 881
rect 1399 884 1404 889
rect 1398 874 1403 879
rect 1426 876 1431 881
rect 1470 876 1475 881
rect 1367 776 1372 781
rect 1397 784 1402 789
rect 1396 774 1401 779
rect 1424 776 1429 781
rect 1468 776 1473 781
rect 1158 724 1163 729
rect 500 674 505 679
rect 530 682 535 687
rect 529 672 534 677
rect 557 674 562 679
rect 601 674 606 679
rect 511 560 516 565
rect 541 568 546 573
rect 540 558 545 563
rect 568 560 573 565
rect 612 560 617 565
rect 1158 670 1163 675
rect 1366 669 1371 674
rect 1396 677 1401 682
rect 1395 667 1400 672
rect 1423 669 1428 674
rect 1467 669 1472 674
rect 1161 600 1166 605
rect 1161 546 1166 551
rect 1366 565 1371 570
rect 1396 573 1401 578
rect 1395 563 1400 568
rect 1423 565 1428 570
rect 1467 565 1472 570
rect 503 451 508 456
rect 533 459 538 464
rect 532 449 537 454
rect 560 451 565 456
rect 604 451 609 456
rect 1155 452 1160 457
rect 1366 450 1371 455
rect 1396 458 1401 463
rect 1395 448 1400 453
rect 1423 450 1428 455
rect 1467 450 1472 455
rect 1155 398 1160 403
rect 508 326 513 331
rect 538 334 543 339
rect 537 324 542 329
rect 565 326 570 331
rect 609 326 614 331
rect 524 215 529 220
rect 554 223 559 228
rect 553 213 558 218
rect 581 215 586 220
rect 625 215 630 220
rect 514 97 519 102
rect 544 105 549 110
rect 543 95 548 100
rect 571 97 576 102
rect 615 97 620 102
<< pm12contact >>
rect 854 1067 859 1072
rect 863 1066 868 1071
rect 994 1067 999 1072
rect 1003 1066 1008 1071
rect 1129 1067 1134 1072
rect 1138 1066 1143 1071
rect 1267 1066 1272 1071
rect 1276 1065 1281 1070
rect 1216 940 1221 945
rect 1225 939 1230 944
rect 1214 707 1219 712
rect 1223 706 1228 711
rect 1217 583 1222 588
rect 1226 582 1231 587
rect 1211 435 1216 440
rect 1220 434 1225 439
<< metal2 >>
rect 799 1078 802 1084
rect 939 1078 942 1084
rect 1074 1078 1077 1084
rect 799 1075 836 1078
rect 939 1075 976 1078
rect 1074 1075 1111 1078
rect 833 1072 836 1075
rect 973 1072 976 1075
rect 1108 1072 1111 1075
rect 1212 1077 1215 1083
rect 1212 1074 1249 1077
rect 833 1069 854 1072
rect 863 1056 866 1066
rect 973 1069 994 1072
rect 1003 1056 1006 1066
rect 1108 1069 1129 1072
rect 1246 1071 1249 1074
rect 1138 1056 1141 1066
rect 1246 1068 1267 1071
rect 800 1053 866 1056
rect 940 1053 1006 1056
rect 1075 1053 1141 1056
rect 1276 1055 1279 1065
rect 800 1035 803 1053
rect 940 1035 943 1053
rect 1075 1035 1078 1053
rect 514 1028 545 1031
rect 1213 1052 1279 1055
rect 1213 1034 1216 1052
rect 514 983 518 1028
rect 541 975 545 1028
rect 463 970 484 974
rect 475 946 481 970
rect 514 946 518 968
rect 585 946 590 970
rect 1161 951 1164 957
rect 1161 948 1198 951
rect 475 943 594 946
rect 1195 945 1198 948
rect 1195 942 1216 945
rect 518 930 549 933
rect 518 885 522 930
rect 545 877 549 930
rect 1225 929 1228 939
rect 1162 926 1228 929
rect 1399 934 1430 937
rect 1162 908 1165 926
rect 1399 889 1403 934
rect 1426 881 1430 934
rect 467 872 488 876
rect 479 848 485 872
rect 1348 876 1369 880
rect 518 848 522 870
rect 589 848 594 872
rect 1360 852 1366 876
rect 1399 852 1403 874
rect 1470 852 1475 876
rect 1360 849 1479 852
rect 479 845 598 848
rect 523 832 554 835
rect 523 787 527 832
rect 550 779 554 832
rect 1397 834 1428 837
rect 1397 789 1401 834
rect 1424 781 1428 834
rect 472 774 493 778
rect 484 750 490 774
rect 1346 776 1367 780
rect 523 750 527 772
rect 594 750 599 774
rect 1358 752 1364 776
rect 1397 752 1401 774
rect 1468 752 1473 776
rect 484 747 603 750
rect 1358 749 1477 752
rect 530 732 561 735
rect 530 687 534 732
rect 557 679 561 732
rect 1396 727 1427 730
rect 1159 718 1162 724
rect 1159 715 1196 718
rect 1193 712 1196 715
rect 1193 709 1214 712
rect 1223 696 1226 706
rect 1160 693 1226 696
rect 479 674 500 678
rect 491 650 497 674
rect 1160 675 1163 693
rect 1396 682 1400 727
rect 530 650 534 672
rect 601 650 606 674
rect 1423 674 1427 727
rect 1345 669 1366 673
rect 491 647 610 650
rect 1357 645 1363 669
rect 1396 645 1400 667
rect 1467 645 1472 669
rect 1357 642 1476 645
rect 1396 623 1427 626
rect 541 618 572 621
rect 541 573 545 618
rect 568 565 572 618
rect 1162 594 1165 600
rect 1162 591 1199 594
rect 1196 588 1199 591
rect 1196 585 1217 588
rect 1226 572 1229 582
rect 1396 578 1400 623
rect 1163 569 1229 572
rect 1423 570 1427 623
rect 490 560 511 564
rect 502 536 508 560
rect 541 536 545 558
rect 612 536 617 560
rect 1163 551 1166 569
rect 1345 565 1366 569
rect 1357 541 1363 565
rect 1396 541 1400 563
rect 1467 541 1472 565
rect 1357 538 1476 541
rect 502 533 621 536
rect 533 509 564 512
rect 533 464 537 509
rect 560 456 564 509
rect 1396 508 1427 511
rect 1396 463 1400 508
rect 482 451 503 455
rect 494 427 500 451
rect 1423 455 1427 508
rect 533 427 537 449
rect 604 427 609 451
rect 1156 446 1159 452
rect 1345 450 1366 454
rect 1156 443 1193 446
rect 1190 440 1193 443
rect 1190 437 1211 440
rect 494 424 613 427
rect 1220 424 1223 434
rect 1157 421 1223 424
rect 1357 426 1363 450
rect 1396 426 1400 448
rect 1467 426 1472 450
rect 1357 423 1476 426
rect 1157 403 1160 421
rect 538 384 569 387
rect 538 339 542 384
rect 565 331 569 384
rect 487 326 508 330
rect 499 302 505 326
rect 538 302 542 324
rect 609 302 614 326
rect 499 299 618 302
rect 554 273 585 276
rect 554 228 558 273
rect 581 220 585 273
rect 503 215 524 219
rect 515 191 521 215
rect 554 191 558 213
rect 625 191 630 215
rect 515 188 634 191
rect 544 155 575 158
rect 544 110 548 155
rect 571 102 575 155
rect 493 97 514 101
rect 505 73 511 97
rect 544 73 548 95
rect 615 73 620 97
rect 505 70 624 73
<< m123contact >>
rect 806 1115 811 1120
rect 946 1115 951 1120
rect 1081 1115 1086 1120
rect 1219 1114 1224 1119
rect 806 1062 811 1067
rect 824 1066 829 1071
rect 946 1062 951 1067
rect 964 1066 969 1071
rect 1081 1062 1086 1067
rect 1099 1066 1104 1071
rect 1219 1061 1224 1066
rect 1237 1065 1242 1070
rect 838 1021 843 1026
rect 978 1021 983 1026
rect 1113 1021 1118 1026
rect 1251 1020 1256 1025
rect 1168 988 1173 993
rect 1168 935 1173 940
rect 1186 939 1191 944
rect 1200 894 1205 899
rect 1166 755 1171 760
rect 1166 702 1171 707
rect 1184 706 1189 711
rect 1198 661 1203 666
rect 1169 631 1174 636
rect 1169 578 1174 583
rect 1187 582 1192 587
rect 1201 537 1206 542
rect 1163 483 1168 488
rect 1163 430 1168 435
rect 1181 434 1186 439
rect 1195 389 1200 394
<< metal3 >>
rect 806 1067 809 1115
rect 829 1066 841 1069
rect 838 1026 841 1066
rect 946 1067 949 1115
rect 969 1066 981 1069
rect 978 1026 981 1066
rect 1081 1067 1084 1115
rect 1104 1066 1116 1069
rect 1113 1026 1116 1066
rect 1219 1066 1222 1114
rect 1242 1065 1254 1068
rect 1251 1025 1254 1065
rect 1168 940 1171 988
rect 1191 939 1203 942
rect 1200 899 1203 939
rect 1166 707 1169 755
rect 1189 706 1201 709
rect 1198 666 1201 706
rect 1169 583 1172 631
rect 1192 582 1204 585
rect 1201 542 1204 582
rect 1163 435 1166 483
rect 1186 434 1198 437
rect 1195 394 1198 434
<< labels >>
rlabel metal1 824 1015 828 1018 1 gnd
rlabel metal1 874 1021 877 1023 1 gnd
rlabel metal1 822 1071 823 1073 1 gnd
rlabel metal1 818 1115 821 1117 5 vdd
rlabel metal1 819 1061 822 1063 1 vdd
rlabel metal1 903 1050 907 1054 7 p0
rlabel metal1 795 1085 796 1088 1 a0
rlabel metal1 795 1031 796 1034 1 b0
rlabel metal1 964 1015 968 1018 1 gnd
rlabel metal1 1014 1021 1017 1023 1 gnd
rlabel metal1 962 1071 963 1073 1 gnd
rlabel metal1 958 1115 961 1117 5 vdd
rlabel metal1 959 1061 962 1063 1 vdd
rlabel metal1 1099 1015 1103 1018 1 gnd
rlabel metal1 1149 1021 1152 1023 1 gnd
rlabel metal1 1097 1071 1098 1073 1 gnd
rlabel metal1 1093 1115 1096 1117 5 vdd
rlabel metal1 1094 1061 1097 1063 1 vdd
rlabel metal1 1237 1014 1241 1017 1 gnd
rlabel metal1 1287 1020 1290 1022 1 gnd
rlabel metal1 1235 1070 1236 1072 1 gnd
rlabel metal1 1231 1114 1234 1116 5 vdd
rlabel metal1 1232 1060 1235 1062 1 vdd
rlabel metal1 935 1031 936 1034 1 b1
rlabel metal1 935 1085 936 1088 1 a1
rlabel metal1 1070 1085 1071 1088 1 a2
rlabel metal1 1070 1031 1071 1034 1 b2
rlabel metal1 1208 1084 1209 1087 1 a3
rlabel metal1 1208 1030 1209 1033 1 b3
rlabel metal1 1316 1049 1320 1053 7 p3
rlabel metal1 1043 1050 1047 1054 1 p1
rlabel metal1 1178 1050 1182 1054 1 p2
rlabel metal1 797 960 798 961 7 g0
rlabel metal1 734 954 735 955 3 b0
rlabel metal1 732 961 733 962 3 a0
rlabel metal1 757 928 757 928 1 gnd!
rlabel metal1 757 992 757 992 5 vdd!
rlabel metal1 797 886 798 887 7 g1
rlabel metal1 757 785 757 785 1 gnd!
rlabel metal1 757 849 757 849 5 vdd!
rlabel metal1 757 711 757 711 1 gnd!
rlabel metal1 757 775 757 775 5 vdd!
rlabel metal1 732 818 733 819 3 a2
rlabel metal1 734 811 735 812 3 b2
rlabel metal1 733 744 734 745 3 a3
rlabel metal1 734 737 735 738 3 b3
rlabel metal1 797 743 798 744 7 g3
rlabel metal1 734 880 735 881 3 b1
rlabel metal1 733 887 734 888 3 a1
rlabel metal1 757 918 757 918 5 vdd!
rlabel metal1 757 854 757 854 1 gnd!
rlabel metal1 1186 888 1190 891 1 gnd
rlabel metal1 1236 894 1239 896 1 gnd
rlabel metal1 1184 944 1185 946 1 gnd
rlabel metal1 1180 988 1183 990 5 vdd
rlabel metal1 1181 934 1184 936 1 vdd
rlabel metal1 1157 958 1158 961 1 p0
rlabel metal1 1157 904 1158 907 1 cin
rlabel metal1 797 817 798 818 7 g2
rlabel metal1 994 898 995 899 1 p3
rlabel metal1 971 898 972 899 1 p2
rlabel metal1 944 898 945 899 1 p1
rlabel metal1 911 898 912 899 1 cin
rlabel metal1 977 821 978 822 1 g3
rlabel metal1 959 820 960 821 1 g2
rlabel metal1 942 820 943 821 1 g1
rlabel metal1 921 820 922 821 1 g0
rlabel metal1 1010 764 1012 765 1 gnd
rlabel metal1 1018 829 1020 830 1 vdd
rlabel metal1 932 898 933 900 1 p0
rlabel metal1 1076 850 1083 851 1 vdd
rlabel metal1 1039 908 1046 909 1 vdd
rlabel metal1 1004 978 1006 979 1 vdd
rlabel metal1 996 913 998 914 1 gnd
rlabel metal1 1026 846 1032 850 1 clk
rlabel metal1 1041 789 1044 822 1 c3
rlabel metal1 1003 896 1014 900 1 c3bar
rlabel metal1 896 819 899 823 3 clk
rlabel metal1 906 816 910 825 1 gnd
rlabel metal1 996 937 1004 941 1 clk_org
rlabel metal1 1012 938 1024 941 1 clk
rlabel metal1 1006 526 1008 527 1 gnd
rlabel metal1 1014 591 1016 592 1 vdd
rlabel metal1 1072 612 1079 613 1 vdd
rlabel metal1 1035 670 1042 671 1 vdd
rlabel metal1 1000 740 1002 741 1 vdd
rlabel metal1 992 675 994 676 1 gnd
rlabel metal1 1022 608 1028 612 1 clk
rlabel metal1 992 699 1000 703 1 clk_org
rlabel metal1 1008 700 1020 703 1 clk
rlabel metal1 984 660 985 661 1 p2
rlabel metal1 957 660 958 661 1 p1
rlabel metal1 924 660 925 661 1 cin
rlabel metal1 972 582 973 583 1 g2
rlabel metal1 955 582 956 583 1 g1
rlabel metal1 934 582 935 583 1 g0
rlabel metal1 945 660 946 662 1 p0
rlabel metal1 909 581 912 585 3 clk
rlabel metal1 919 578 923 587 1 gnd
rlabel metal1 1011 299 1013 300 1 gnd
rlabel metal1 1019 364 1021 365 1 vdd
rlabel metal1 1077 385 1084 386 1 vdd
rlabel metal1 1040 443 1047 444 1 vdd
rlabel metal1 1005 513 1007 514 1 vdd
rlabel metal1 997 448 999 449 1 gnd
rlabel metal1 1027 381 1033 385 1 clk
rlabel metal1 997 472 1005 476 1 clk_org
rlabel metal1 1013 473 1025 476 1 clk
rlabel metal1 998 550 1002 614 1 c2bar
rlabel metal1 1037 551 1040 584 1 c2
rlabel metal1 951 351 955 360 1 gnd
rlabel metal1 941 354 944 358 3 clk
rlabel metal1 977 433 978 435 1 p0
rlabel metal1 966 355 967 356 1 g0
rlabel metal1 987 355 988 356 1 g1
rlabel metal1 956 433 957 434 1 cin
rlabel metal1 989 433 990 434 1 p1
rlabel metal1 1002 371 1009 378 1 c1bar
rlabel metal1 1042 324 1045 357 1 c1
rlabel metal1 1013 76 1015 77 1 gnd
rlabel metal1 1021 141 1023 142 1 vdd
rlabel metal1 1079 162 1086 163 1 vdd
rlabel metal1 1042 220 1049 221 1 vdd
rlabel metal1 1007 290 1009 291 1 vdd
rlabel metal1 999 225 1001 226 1 gnd
rlabel metal1 1029 158 1035 162 1 clk
rlabel metal1 999 249 1007 253 1 clk_org
rlabel metal1 1015 250 1027 253 1 clk
rlabel metal1 972 128 976 137 1 gnd
rlabel metal1 962 131 965 135 3 clk
rlabel metal1 998 210 999 212 1 p0
rlabel metal1 987 132 988 133 1 g0
rlabel metal1 977 210 978 211 1 cin
rlabel metal1 996 151 1053 155 1 c0bar
rlabel metal1 1044 101 1047 134 1 c0
rlabel metal2 480 971 480 971 1 clk_org
rlabel metal1 499 1022 501 1023 5 vdd
rlabel metal1 493 950 496 951 1 gnd
rlabel metal2 484 873 484 873 1 clk_org
rlabel metal1 503 924 505 925 5 vdd
rlabel metal1 497 852 500 853 1 gnd
rlabel metal2 489 775 489 775 1 clk_org
rlabel metal1 508 826 510 827 5 vdd
rlabel metal1 502 754 505 755 1 gnd
rlabel metal2 496 675 496 675 1 clk_org
rlabel metal1 515 726 517 727 5 vdd
rlabel metal1 509 654 512 655 1 gnd
rlabel metal1 520 540 523 541 1 gnd
rlabel metal1 526 612 528 613 5 vdd
rlabel metal2 507 561 507 561 1 clk_org
rlabel metal1 512 431 515 432 1 gnd
rlabel metal1 518 503 520 504 5 vdd
rlabel metal2 499 452 499 452 1 clk_org
rlabel metal1 517 306 520 307 1 gnd
rlabel metal1 523 378 525 379 5 vdd
rlabel metal2 504 327 504 327 1 clk_org
rlabel metal1 533 195 536 196 1 gnd
rlabel metal1 539 267 541 268 5 vdd
rlabel metal2 520 216 520 216 1 clk_org
rlabel metal1 523 77 526 78 1 gnd
rlabel metal1 529 149 531 150 5 vdd
rlabel metal2 510 98 510 98 1 clk_org
rlabel metal1 1378 856 1381 857 1 gnd
rlabel metal1 1384 928 1386 929 5 vdd
rlabel metal2 1365 877 1365 877 1 clk_org
rlabel metal1 479 980 479 980 1 cinin
rlabel metal1 633 977 633 977 1 cin
rlabel metal1 487 882 487 882 1 a0in
rlabel metal1 636 879 636 879 1 a0
rlabel metal1 490 784 490 784 1 b0in
rlabel metal1 643 781 643 781 1 b0
rlabel metal1 498 685 498 685 1 a1in
rlabel metal1 649 680 649 680 1 a1
rlabel metal1 509 570 509 570 1 b1in
rlabel metal1 662 567 662 567 1 b1
rlabel metal1 501 462 501 462 1 a2in
rlabel metal1 652 458 652 458 1 a2
rlabel metal1 506 336 506 336 1 b2in
rlabel metal1 658 333 658 333 1 b2
rlabel metal1 521 225 521 225 1 a3in
rlabel metal1 675 221 675 221 1 a3
rlabel metal1 513 106 513 106 1 b3in
rlabel metal1 664 105 664 105 1 b3
rlabel metal1 1365 885 1365 885 1 s0in
rlabel metal1 1376 756 1379 757 1 gnd
rlabel metal1 1382 828 1384 829 5 vdd
rlabel metal2 1363 777 1363 777 1 clk_org
rlabel metal1 1375 649 1378 650 1 gnd
rlabel metal1 1381 721 1383 722 5 vdd
rlabel metal2 1362 670 1362 670 1 clk_org
rlabel metal1 1375 545 1378 546 1 gnd
rlabel metal1 1381 617 1383 618 5 vdd
rlabel metal2 1362 566 1362 566 1 clk_org
rlabel metal1 1375 430 1378 431 1 gnd
rlabel metal1 1381 502 1383 503 5 vdd
rlabel metal2 1362 451 1362 451 1 clk_org
rlabel metal1 1187 531 1191 534 1 gnd
rlabel metal1 1237 537 1240 539 1 gnd
rlabel metal1 1185 587 1186 589 1 gnd
rlabel metal1 1181 631 1184 633 5 vdd
rlabel metal1 1182 577 1185 579 1 vdd
rlabel metal1 1158 601 1159 604 1 p2
rlabel metal1 1158 547 1159 550 1 c1
rlabel metal1 1152 399 1153 402 1 c0
rlabel metal1 1179 439 1180 441 1 gnd
rlabel metal1 1152 453 1153 456 1 p1
rlabel metal1 1176 429 1179 431 1 vdd
rlabel metal1 1175 483 1178 485 5 vdd
rlabel metal1 1231 389 1234 391 1 gnd
rlabel metal1 1181 383 1185 386 1 gnd
rlabel metal1 1155 725 1156 728 1 p3
rlabel metal1 1155 671 1156 674 1 c2
rlabel metal1 1179 701 1182 703 1 vdd
rlabel metal1 1178 755 1181 757 5 vdd
rlabel metal1 1182 711 1183 713 1 gnd
rlabel metal1 1234 661 1237 663 1 gnd
rlabel metal1 1184 655 1188 658 1 gnd
rlabel metal1 1515 881 1515 881 1 s0
rlabel metal1 1364 786 1364 786 1 c3
rlabel metal1 1517 782 1517 782 7 cout
rlabel metal1 1363 678 1363 678 1 s3in
rlabel metal1 1516 675 1516 675 1 s3
rlabel metal1 1363 575 1363 575 1 s2in
rlabel metal1 1515 572 1515 572 1 s2
rlabel metal1 1365 459 1365 459 1 s1in
rlabel metal1 1516 456 1516 456 1 s1
rlabel metal1 1268 420 1268 420 1 s1in
rlabel metal1 1274 568 1274 568 1 s2in
rlabel metal1 1273 692 1273 692 1 s3in
rlabel metal1 1586 823 1588 824 1 vdd
rlabel metal1 1578 758 1580 759 1 gnd
rlabel metal1 1588 724 1590 725 1 vdd
rlabel metal1 1580 659 1582 660 1 gnd
rlabel metal1 1584 622 1586 623 1 vdd
rlabel metal1 1576 557 1578 558 1 gnd
rlabel metal1 1581 503 1583 504 1 vdd
rlabel metal1 1573 438 1575 439 1 gnd
rlabel metal1 1582 926 1584 927 1 vdd
rlabel metal1 1574 861 1576 862 1 gnd
rlabel metal1 1579 582 1579 582 1 s2
rlabel metal1 1577 463 1577 463 1 s1
rlabel metal1 1587 684 1587 684 1 s3
rlabel metal1 1581 783 1581 783 1 cout
rlabel metal1 1579 888 1579 888 1 s0
rlabel metal1 1269 925 1269 925 1 s0in
<< end >>
